//*******************************************************************************
// Project      : 
// Module       : div2.v
// Description  : frequency divider - 2 
// Designer     :
// Version      : 
//********************************************************************************

module div2(
input		in,
output		out
);

wire d0;
//*********************************************************************
//
// D flip flop
//
//*********************************************************************
FFDHD2X u0(.CK(in), .D(d0), .Q(out), .QN(d0));


//********************************************************************************
//
// END of Module
//
//********************************************************************************
endmodule
