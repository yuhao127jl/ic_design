
//----------------------------------------------------------//
//
// include file
//
//----------------------------------------------------------//






//----------------------------------------------------------//
//
// router env
//
//----------------------------------------------------------//
class router_env extends uvm_env;




endclass






