
typedef uvm_sequencer #(packet_transaction) packet_sequencer;

