//*******************************************************************************
// Project		: 
// Module		: cos_tbl.v
// Description	: 
// Designer		: 
// Version		: 
//*******************************************************************************

module cos_tbl(
    input wire[9:0]      addr,
    output reg[15:0]     cos_dat
);

//**********************************************************
//
// always
//
//**********************************************************
always @(*)
begin
    case(addr)
    10'd0       : cos_dat = 16'b0111111110100110;  
    10'd1       : cos_dat = 16'b0111111110100101;  
    10'd2       : cos_dat = 16'b0111111110100011;  
    10'd3       : cos_dat = 16'b0111111110100000;  
    10'd4       : cos_dat = 16'b0111111110011100;  
    10'd5       : cos_dat = 16'b0111111110010110;  
    10'd6       : cos_dat = 16'b0111111110001111;  
    10'd7       : cos_dat = 16'b0111111110000111;  
    10'd8       : cos_dat = 16'b0111111101111110;  
    10'd9       : cos_dat = 16'b0111111101110100;  
    10'd10      : cos_dat = 16'b0111111101101000;  
    10'd11      : cos_dat = 16'b0111111101011011;  
    10'd12      : cos_dat = 16'b0111111101001101;  
    10'd13      : cos_dat = 16'b0111111100111101;  
    10'd14      : cos_dat = 16'b0111111100101101;  
    10'd15      : cos_dat = 16'b0111111100011011;  
    10'd16      : cos_dat = 16'b0111111100001000;  
    10'd17      : cos_dat = 16'b0111111011110100;  
    10'd18      : cos_dat = 16'b0111111011011110;  
    10'd19      : cos_dat = 16'b0111111011000111;  
    10'd20      : cos_dat = 16'b0111111010110000;  
    10'd21      : cos_dat = 16'b0111111010010110;  
    10'd22      : cos_dat = 16'b0111111001111100;  
    10'd23      : cos_dat = 16'b0111111001100000;  
    10'd24      : cos_dat = 16'b0111111001000011;  
    10'd25      : cos_dat = 16'b0111111000100101;  
    10'd26      : cos_dat = 16'b0111111000000110;  
    10'd27      : cos_dat = 16'b0111110111100110;  
    10'd28      : cos_dat = 16'b0111110111000100;  
    10'd29      : cos_dat = 16'b0111110110100001;  
    10'd30      : cos_dat = 16'b0111110101111101;  
    10'd31      : cos_dat = 16'b0111110101011000;  
    10'd32      : cos_dat = 16'b0111110100110001;  
    10'd33      : cos_dat = 16'b0111110100001001;  
    10'd34      : cos_dat = 16'b0111110011100000;  
    10'd35      : cos_dat = 16'b0111110010110110;  
    10'd36      : cos_dat = 16'b0111110010001011;  
    10'd37      : cos_dat = 16'b0111110001011110;  
    10'd38      : cos_dat = 16'b0111110000110000;  
    10'd39      : cos_dat = 16'b0111110000000001;  
    10'd40      : cos_dat = 16'b0111101111010001;  
    10'd41      : cos_dat = 16'b0111101110100000;  
    10'd42      : cos_dat = 16'b0111101101101101;  
    10'd43      : cos_dat = 16'b0111101100111010;  
    10'd44      : cos_dat = 16'b0111101100000101;  
    10'd45      : cos_dat = 16'b0111101011001111;  
    10'd46      : cos_dat = 16'b0111101010010111;  
    10'd47      : cos_dat = 16'b0111101001011111;  
    10'd48      : cos_dat = 16'b0111101000100101;  
    10'd49      : cos_dat = 16'b0111100111101010;  
    10'd50      : cos_dat = 16'b0111100110101110;  
    10'd51      : cos_dat = 16'b0111100101110001;  
    10'd52      : cos_dat = 16'b0111100100110011;  
    10'd53      : cos_dat = 16'b0111100011110011;  
    10'd54      : cos_dat = 16'b0111100010110010;  
    10'd55      : cos_dat = 16'b0111100001110001;  
    10'd56      : cos_dat = 16'b0111100000101101;  
    10'd57      : cos_dat = 16'b0111011111101001;  
    10'd58      : cos_dat = 16'b0111011110100100;  
    10'd59      : cos_dat = 16'b0111011101011101;  
    10'd60      : cos_dat = 16'b0111011100010110;  
    10'd61      : cos_dat = 16'b0111011011001101;  
    10'd62      : cos_dat = 16'b0111011010000011;  
    10'd63      : cos_dat = 16'b0111011000111000;  
    10'd64      : cos_dat = 16'b0111010111101100;  
    10'd65      : cos_dat = 16'b0111010110011110;  
    10'd66      : cos_dat = 16'b0111010101010000;  
    10'd67      : cos_dat = 16'b0111010100000000;  
    10'd68      : cos_dat = 16'b0111010010101111;  
    10'd69      : cos_dat = 16'b0111010001011110;  
    10'd70      : cos_dat = 16'b0111010000001011;  
    10'd71      : cos_dat = 16'b0111001110110110;  
    10'd72      : cos_dat = 16'b0111001101100001;  
    10'd73      : cos_dat = 16'b0111001100001011;  
    10'd74      : cos_dat = 16'b0111001010110011;  
    10'd75      : cos_dat = 16'b0111001001011011;  
    10'd76      : cos_dat = 16'b0111001000000001;  
    10'd77      : cos_dat = 16'b0111000110100110;  
    10'd78      : cos_dat = 16'b0111000101001010;  
    10'd79      : cos_dat = 16'b0111000011101101;  
    10'd80      : cos_dat = 16'b0111000010001111;  
    10'd81      : cos_dat = 16'b0111000000110000;  
    10'd82      : cos_dat = 16'b0110111111010000;  
    10'd83      : cos_dat = 16'b0110111101101111;  
    10'd84      : cos_dat = 16'b0110111100001100;  
    10'd85      : cos_dat = 16'b0110111010101001;  
    10'd86      : cos_dat = 16'b0110111001000100;  
    10'd87      : cos_dat = 16'b0110110111011111;  
    10'd88      : cos_dat = 16'b0110110101111000;  
    10'd89      : cos_dat = 16'b0110110100010000;  
    10'd90      : cos_dat = 16'b0110110010101000;  
    10'd91      : cos_dat = 16'b0110110000111110;  
    10'd92      : cos_dat = 16'b0110101111010011;  
    10'd93      : cos_dat = 16'b0110101101100111;  
    10'd94      : cos_dat = 16'b0110101011111010;  
    10'd95      : cos_dat = 16'b0110101010001100;  
    10'd96      : cos_dat = 16'b0110101000011101;  
    10'd97      : cos_dat = 16'b0110100110101101;  
    10'd98      : cos_dat = 16'b0110100100111100;  
    10'd99      : cos_dat = 16'b0110100011001010;  
    10'd100     : cos_dat = 16'b0110100001010111;  
    10'd101     : cos_dat = 16'b0110011111100011;  
    10'd102     : cos_dat = 16'b0110011101101110;  
    10'd103     : cos_dat = 16'b0110011011111000;  
    10'd104     : cos_dat = 16'b0110011010000001;  
    10'd105     : cos_dat = 16'b0110011000001001;  
    10'd106     : cos_dat = 16'b0110010110010000;  
    10'd107     : cos_dat = 16'b0110010100010110;  
    10'd108     : cos_dat = 16'b0110010010011011;  
    10'd109     : cos_dat = 16'b0110010000011111;  
    10'd110     : cos_dat = 16'b0110001110100010;  
    10'd111     : cos_dat = 16'b0110001100100100;  
    10'd112     : cos_dat = 16'b0110001010100101;  
    10'd113     : cos_dat = 16'b0110001000100101;  
    10'd114     : cos_dat = 16'b0110000110100101;  
    10'd115     : cos_dat = 16'b0110000100100011;  
    10'd116     : cos_dat = 16'b0110000010100000;  
    10'd117     : cos_dat = 16'b0110000000011101;  
    10'd118     : cos_dat = 16'b0101111110011000;  
    10'd119     : cos_dat = 16'b0101111100010011;  
    10'd120     : cos_dat = 16'b0101111010001101;  
    10'd121     : cos_dat = 16'b0101111000000101;  
    10'd122     : cos_dat = 16'b0101110101111101;  
    10'd123     : cos_dat = 16'b0101110011110100;  
    10'd124     : cos_dat = 16'b0101110001101010;  
    10'd125     : cos_dat = 16'b0101101111100000;  
    10'd126     : cos_dat = 16'b0101101101010100;  
    10'd127     : cos_dat = 16'b0101101011000111;  
    10'd128     : cos_dat = 16'b0101101000111010;  
    10'd129     : cos_dat = 16'b0101100110101011;  
    10'd130     : cos_dat = 16'b0101100100011100;  
    10'd131     : cos_dat = 16'b0101100010001100;  
    10'd132     : cos_dat = 16'b0101011111111011;  
    10'd133     : cos_dat = 16'b0101011101101010;  
    10'd134     : cos_dat = 16'b0101011011010111;  
    10'd135     : cos_dat = 16'b0101011001000011;  
    10'd136     : cos_dat = 16'b0101010110101111;  
    10'd137     : cos_dat = 16'b0101010100011010;  
    10'd138     : cos_dat = 16'b0101010010000100;  
    10'd139     : cos_dat = 16'b0101001111101101;  
    10'd140     : cos_dat = 16'b0101001101010110;  
    10'd141     : cos_dat = 16'b0101001010111110;  
    10'd142     : cos_dat = 16'b0101001000100100;  
    10'd143     : cos_dat = 16'b0101000110001010;  
    10'd144     : cos_dat = 16'b0101000011110000;  
    10'd145     : cos_dat = 16'b0101000001010100;  
    10'd146     : cos_dat = 16'b0100111110111000;  
    10'd147     : cos_dat = 16'b0100111100011011;  
    10'd148     : cos_dat = 16'b0100111001111101;  
    10'd149     : cos_dat = 16'b0100110111011110;  
    10'd150     : cos_dat = 16'b0100110100111111;  
    10'd151     : cos_dat = 16'b0100110010011111;  
    10'd152     : cos_dat = 16'b0100101111111110;  
    10'd153     : cos_dat = 16'b0100101101011101;  
    10'd154     : cos_dat = 16'b0100101010111010;  
    10'd155     : cos_dat = 16'b0100101000010111;  
    10'd156     : cos_dat = 16'b0100100101110100;  
    10'd157     : cos_dat = 16'b0100100011001111;  
    10'd158     : cos_dat = 16'b0100100000101010;  
    10'd159     : cos_dat = 16'b0100011110000100;  
    10'd160     : cos_dat = 16'b0100011011011110;  
    10'd161     : cos_dat = 16'b0100011000110111;  
    10'd162     : cos_dat = 16'b0100010110001111;  
    10'd163     : cos_dat = 16'b0100010011100110;  
    10'd164     : cos_dat = 16'b0100010000111101;  
    10'd165     : cos_dat = 16'b0100001110010011;  
    10'd166     : cos_dat = 16'b0100001011101001;  
    10'd167     : cos_dat = 16'b0100001000111110;  
    10'd168     : cos_dat = 16'b0100000110010010;  
    10'd169     : cos_dat = 16'b0100000011100101;  
    10'd170     : cos_dat = 16'b0100000000111000;  
    10'd171     : cos_dat = 16'b0011111110001011;  
    10'd172     : cos_dat = 16'b0011111011011100;  
    10'd173     : cos_dat = 16'b0011111000101101;  
    10'd174     : cos_dat = 16'b0011110101111110;  
    10'd175     : cos_dat = 16'b0011110011001110;  
    10'd176     : cos_dat = 16'b0011110000011101;  
    10'd177     : cos_dat = 16'b0011101101101100;  
    10'd178     : cos_dat = 16'b0011101010111010;  
    10'd179     : cos_dat = 16'b0011101000001000;  
    10'd180     : cos_dat = 16'b0011100101010101;  
    10'd181     : cos_dat = 16'b0011100010100001;  
    10'd182     : cos_dat = 16'b0011011111101101;  
    10'd183     : cos_dat = 16'b0011011100111001;  
    10'd184     : cos_dat = 16'b0011011010000011;  
    10'd185     : cos_dat = 16'b0011010111001110;  
    10'd186     : cos_dat = 16'b0011010100011000;  
    10'd187     : cos_dat = 16'b0011010001100001;  
    10'd188     : cos_dat = 16'b0011001110101010;  
    10'd189     : cos_dat = 16'b0011001011110010;  
    10'd190     : cos_dat = 16'b0011001000111010;  
    10'd191     : cos_dat = 16'b0011000110000001;  
    10'd192     : cos_dat = 16'b0011000011001000;  
    10'd193     : cos_dat = 16'b0011000000001110;  
    10'd194     : cos_dat = 16'b0010111101010100;  
    10'd195     : cos_dat = 16'b0010111010011010;  
    10'd196     : cos_dat = 16'b0010110111011111;  
    10'd197     : cos_dat = 16'b0010110100100011;  
    10'd198     : cos_dat = 16'b0010110001101000;  
    10'd199     : cos_dat = 16'b0010101110101011;  
    10'd200     : cos_dat = 16'b0010101011101111;  
    10'd201     : cos_dat = 16'b0010101000110010;  
    10'd202     : cos_dat = 16'b0010100101110100;  
    10'd203     : cos_dat = 16'b0010100010110110;  
    10'd204     : cos_dat = 16'b0010011111111000;  
    10'd205     : cos_dat = 16'b0010011100111001;  
    10'd206     : cos_dat = 16'b0010011001111010;  
    10'd207     : cos_dat = 16'b0010010110111010;  
    10'd208     : cos_dat = 16'b0010010011111011;  
    10'd209     : cos_dat = 16'b0010010000111010;  
    10'd210     : cos_dat = 16'b0010001101111010;  
    10'd211     : cos_dat = 16'b0010001010111001;  
    10'd212     : cos_dat = 16'b0010000111111000;  
    10'd213     : cos_dat = 16'b0010000100110110;  
    10'd214     : cos_dat = 16'b0010000001110100;  
    10'd215     : cos_dat = 16'b0001111110110010;  
    10'd216     : cos_dat = 16'b0001111011110000;  
    10'd217     : cos_dat = 16'b0001111000101101;  
    10'd218     : cos_dat = 16'b0001110101101010;  
    10'd219     : cos_dat = 16'b0001110010100111;  
    10'd220     : cos_dat = 16'b0001101111100011;  
    10'd221     : cos_dat = 16'b0001101100011111;  
    10'd222     : cos_dat = 16'b0001101001011011;  
    10'd223     : cos_dat = 16'b0001100110010111;  
    10'd224     : cos_dat = 16'b0001100011010010;  
    10'd225     : cos_dat = 16'b0001100000001101;  
    10'd226     : cos_dat = 16'b0001011101001000;  
    10'd227     : cos_dat = 16'b0001011010000011;  
    10'd228     : cos_dat = 16'b0001010110111101;  
    10'd229     : cos_dat = 16'b0001010011110111;  
    10'd230     : cos_dat = 16'b0001010000110001;  
    10'd231     : cos_dat = 16'b0001001101101011;  
    10'd232     : cos_dat = 16'b0001001010100101;  
    10'd233     : cos_dat = 16'b0001000111011110;  
    10'd234     : cos_dat = 16'b0001000100010111;  
    10'd235     : cos_dat = 16'b0001000001010001;  
    10'd236     : cos_dat = 16'b0000111110001010;  
    10'd237     : cos_dat = 16'b0000111011000010;  
    10'd238     : cos_dat = 16'b0000110111111011;  
    10'd239     : cos_dat = 16'b0000110100110100;  
    10'd240     : cos_dat = 16'b0000110001101100;  
    10'd241     : cos_dat = 16'b0000101110100100;  
    10'd242     : cos_dat = 16'b0000101011011100;  
    10'd243     : cos_dat = 16'b0000101000010101;  
    10'd244     : cos_dat = 16'b0000100101001101;  
    10'd245     : cos_dat = 16'b0000100010000100;  
    10'd246     : cos_dat = 16'b0000011110111100;  
    10'd247     : cos_dat = 16'b0000011011110100;  
    10'd248     : cos_dat = 16'b0000011000101100;  
    10'd249     : cos_dat = 16'b0000010101100011;  
    10'd250     : cos_dat = 16'b0000010010011011;  
    10'd251     : cos_dat = 16'b0000001111010010;  
    10'd252     : cos_dat = 16'b0000001100001010;  
    10'd253     : cos_dat = 16'b0000001001000001;  
    10'd254     : cos_dat = 16'b0000000101111001;  
    10'd255     : cos_dat = 16'b0000000010110000;  
    10'd256     : cos_dat = 16'b1111111111100111;  
    10'd257     : cos_dat = 16'b1111111100011111;  
    10'd258     : cos_dat = 16'b1111111001010110;  
    10'd259     : cos_dat = 16'b1111110110001110;  
    10'd260     : cos_dat = 16'b1111110011000101;  
    10'd261     : cos_dat = 16'b1111101111111101;  
    10'd262     : cos_dat = 16'b1111101100110100;  
    10'd263     : cos_dat = 16'b1111101001101100;  
    10'd264     : cos_dat = 16'b1111100110100011;  
    10'd265     : cos_dat = 16'b1111100011011011;  
    10'd266     : cos_dat = 16'b1111100000010011;  
    10'd267     : cos_dat = 16'b1111011101001010;  
    10'd268     : cos_dat = 16'b1111011010000010;  
    10'd269     : cos_dat = 16'b1111010110111010;  
    10'd270     : cos_dat = 16'b1111010011110010;  
    10'd271     : cos_dat = 16'b1111010000101011;  
    10'd272     : cos_dat = 16'b1111001101100011;  
    10'd273     : cos_dat = 16'b1111001010011011;  
    10'd274     : cos_dat = 16'b1111000111010100;  
    10'd275     : cos_dat = 16'b1111000100001101;  
    10'd276     : cos_dat = 16'b1111000001000110;  
    10'd277     : cos_dat = 16'b1110111101111111;  
    10'd278     : cos_dat = 16'b1110111010111000;  
    10'd279     : cos_dat = 16'b1110110111110001;  
    10'd280     : cos_dat = 16'b1110110100101011;  
    10'd281     : cos_dat = 16'b1110110001100100;  
    10'd282     : cos_dat = 16'b1110101110011110;  
    10'd283     : cos_dat = 16'b1110101011011000;  
    10'd284     : cos_dat = 16'b1110101000010010;  
    10'd285     : cos_dat = 16'b1110100101001101;  
    10'd286     : cos_dat = 16'b1110100010001000;  
    10'd287     : cos_dat = 16'b1110011111000011;  
    10'd288     : cos_dat = 16'b1110011011111110;  
    10'd289     : cos_dat = 16'b1110011000111001;  
    10'd290     : cos_dat = 16'b1110010101110101;  
    10'd291     : cos_dat = 16'b1110010010110001;  
    10'd292     : cos_dat = 16'b1110001111101101;  
    10'd293     : cos_dat = 16'b1110001100101001;  
    10'd294     : cos_dat = 16'b1110001001100110;  
    10'd295     : cos_dat = 16'b1110000110100011;  
    10'd296     : cos_dat = 16'b1110000011100000;  
    10'd297     : cos_dat = 16'b1110000000011110;  
    10'd298     : cos_dat = 16'b1101111101011100;  
    10'd299     : cos_dat = 16'b1101111010011010;  
    10'd300     : cos_dat = 16'b1101110111011001;  
    10'd301     : cos_dat = 16'b1101110100010111;  
    10'd302     : cos_dat = 16'b1101110001010111;  
    10'd303     : cos_dat = 16'b1101101110010110;  
    10'd304     : cos_dat = 16'b1101101011010110;  
    10'd305     : cos_dat = 16'b1101101000010110;  
    10'd306     : cos_dat = 16'b1101100101010111;  
    10'd307     : cos_dat = 16'b1101100010011000;  
    10'd308     : cos_dat = 16'b1101011111011001;  
    10'd309     : cos_dat = 16'b1101011100011011;  
    10'd310     : cos_dat = 16'b1101011001011101;  
    10'd311     : cos_dat = 16'b1101010110100000;  
    10'd312     : cos_dat = 16'b1101010011100011;  
    10'd313     : cos_dat = 16'b1101010000100110;  
    10'd314     : cos_dat = 16'b1101001101101010;  
    10'd315     : cos_dat = 16'b1101001010101110;  
    10'd316     : cos_dat = 16'b1101000111110011;  
    10'd317     : cos_dat = 16'b1101000100111000;  
    10'd318     : cos_dat = 16'b1101000001111110;  
    10'd319     : cos_dat = 16'b1100111111000100;  
    10'd320     : cos_dat = 16'b1100111100001010;  
    10'd321     : cos_dat = 16'b1100111001010001;  
    10'd322     : cos_dat = 16'b1100110110011001;  
    10'd323     : cos_dat = 16'b1100110011100001;  
    10'd324     : cos_dat = 16'b1100110000101001;  
    10'd325     : cos_dat = 16'b1100101101110010;  
    10'd326     : cos_dat = 16'b1100101010111011;  
    10'd327     : cos_dat = 16'b1100101000000101;  
    10'd328     : cos_dat = 16'b1100100101010000;  
    10'd329     : cos_dat = 16'b1100100010011011;  
    10'd330     : cos_dat = 16'b1100011111100110;  
    10'd331     : cos_dat = 16'b1100011100110011;  
    10'd332     : cos_dat = 16'b1100011001111111;  
    10'd333     : cos_dat = 16'b1100010111001100;  
    10'd334     : cos_dat = 16'b1100010100011010;  
    10'd335     : cos_dat = 16'b1100010001101000;  
    10'd336     : cos_dat = 16'b1100001110110111;  
    10'd337     : cos_dat = 16'b1100001100000111;  
    10'd338     : cos_dat = 16'b1100001001010111;  
    10'd339     : cos_dat = 16'b1100000110100111;  
    10'd340     : cos_dat = 16'b1100000011111001;  
    10'd341     : cos_dat = 16'b1100000001001011;  
    10'd342     : cos_dat = 16'b1011111110011101;  
    10'd343     : cos_dat = 16'b1011111011110000;  
    10'd344     : cos_dat = 16'b1011111001000100;  
    10'd345     : cos_dat = 16'b1011110110011000;  
    10'd346     : cos_dat = 16'b1011110011101101;  
    10'd347     : cos_dat = 16'b1011110001000011;  
    10'd348     : cos_dat = 16'b1011101110011001;  
    10'd349     : cos_dat = 16'b1011101011110000;  
    10'd350     : cos_dat = 16'b1011101001001000;  
    10'd351     : cos_dat = 16'b1011100110100000;  
    10'd352     : cos_dat = 16'b1011100011111001;  
    10'd353     : cos_dat = 16'b1011100001010011;  
    10'd354     : cos_dat = 16'b1011011110101101;  
    10'd355     : cos_dat = 16'b1011011100001000;  
    10'd356     : cos_dat = 16'b1011011001100100;  
    10'd357     : cos_dat = 16'b1011010111000000;  
    10'd358     : cos_dat = 16'b1011010100011101;  
    10'd359     : cos_dat = 16'b1011010001111011;  
    10'd360     : cos_dat = 16'b1011001111011010;  
    10'd361     : cos_dat = 16'b1011001100111001;  
    10'd362     : cos_dat = 16'b1011001010011001;  
    10'd363     : cos_dat = 16'b1011000111111010;  
    10'd364     : cos_dat = 16'b1011000101011100;  
    10'd365     : cos_dat = 16'b1011000010111110;  
    10'd366     : cos_dat = 16'b1011000000100001;  
    10'd367     : cos_dat = 16'b1010111110000101;  
    10'd368     : cos_dat = 16'b1010111011101010;  
    10'd369     : cos_dat = 16'b1010111001001111;  
    10'd370     : cos_dat = 16'b1010110110110110;  
    10'd371     : cos_dat = 16'b1010110100011101;  
    10'd372     : cos_dat = 16'b1010110010000101;  
    10'd373     : cos_dat = 16'b1010101111101101;  
    10'd374     : cos_dat = 16'b1010101101010111;  
    10'd375     : cos_dat = 16'b1010101011000001;  
    10'd376     : cos_dat = 16'b1010101000101100;  
    10'd377     : cos_dat = 16'b1010100110011000;  
    10'd378     : cos_dat = 16'b1010100100000101;  
    10'd379     : cos_dat = 16'b1010100001110010;  
    10'd380     : cos_dat = 16'b1010011111100001;  
    10'd381     : cos_dat = 16'b1010011101010000;  
    10'd382     : cos_dat = 16'b1010011011000000;  
    10'd383     : cos_dat = 16'b1010011000110001;  
    10'd384     : cos_dat = 16'b1010010110100011;  
    10'd385     : cos_dat = 16'b1010010100010110;  
    10'd386     : cos_dat = 16'b1010010010001001;  
    10'd387     : cos_dat = 16'b1010001111111110;  
    10'd388     : cos_dat = 16'b1010001101110011;  
    10'd389     : cos_dat = 16'b1010001011101010;  
    10'd390     : cos_dat = 16'b1010001001100001;  
    10'd391     : cos_dat = 16'b1010000111011001;  
    10'd392     : cos_dat = 16'b1010000101010010;  
    10'd393     : cos_dat = 16'b1010000011001100;  
    10'd394     : cos_dat = 16'b1010000001000111;  
    10'd395     : cos_dat = 16'b1001111111000010;  
    10'd396     : cos_dat = 16'b1001111100111111;  
    10'd397     : cos_dat = 16'b1001111010111101;  
    10'd398     : cos_dat = 16'b1001111000111011;  
    10'd399     : cos_dat = 16'b1001110110111011;  
    10'd400     : cos_dat = 16'b1001110100111011;  
    10'd401     : cos_dat = 16'b1001110010111101;  
    10'd402     : cos_dat = 16'b1001110000111111;  
    10'd403     : cos_dat = 16'b1001101111000010;  
    10'd404     : cos_dat = 16'b1001101101000111;  
    10'd405     : cos_dat = 16'b1001101011001100;  
    10'd406     : cos_dat = 16'b1001101001010010;  
    10'd407     : cos_dat = 16'b1001100111011001;  
    10'd408     : cos_dat = 16'b1001100101100001;  
    10'd409     : cos_dat = 16'b1001100011101011;  
    10'd410     : cos_dat = 16'b1001100001110101;  
    10'd411     : cos_dat = 16'b1001100000000000;  
    10'd412     : cos_dat = 16'b1001011110001100;  
    10'd413     : cos_dat = 16'b1001011100011001;  
    10'd414     : cos_dat = 16'b1001011010101000;  
    10'd415     : cos_dat = 16'b1001011000110111;  
    10'd416     : cos_dat = 16'b1001010111000111;  
    10'd417     : cos_dat = 16'b1001010101011000;  
    10'd418     : cos_dat = 16'b1001010011101011;  
    10'd419     : cos_dat = 16'b1001010001111110;  
    10'd420     : cos_dat = 16'b1001010000010010;  
    10'd421     : cos_dat = 16'b1001001110101000;  
    10'd422     : cos_dat = 16'b1001001100111110;  
    10'd423     : cos_dat = 16'b1001001011010110;  
    10'd424     : cos_dat = 16'b1001001001101110;  
    10'd425     : cos_dat = 16'b1001001000001000;  
    10'd426     : cos_dat = 16'b1001000110100010;  
    10'd427     : cos_dat = 16'b1001000100111110;  
    10'd428     : cos_dat = 16'b1001000011011011;  
    10'd429     : cos_dat = 16'b1001000001111001;  
    10'd430     : cos_dat = 16'b1001000000011000;  
    10'd431     : cos_dat = 16'b1000111110111000;  
    10'd432     : cos_dat = 16'b1000111101011001;  
    10'd433     : cos_dat = 16'b1000111011111011;  
    10'd434     : cos_dat = 16'b1000111010011110;  
    10'd435     : cos_dat = 16'b1000111001000011;  
    10'd436     : cos_dat = 16'b1000110111101000;  
    10'd437     : cos_dat = 16'b1000110110001111;  
    10'd438     : cos_dat = 16'b1000110100110111;  
    10'd439     : cos_dat = 16'b1000110011011111;  
    10'd440     : cos_dat = 16'b1000110010001001;  
    10'd441     : cos_dat = 16'b1000110000110100;  
    10'd442     : cos_dat = 16'b1000101111100000;  
    10'd443     : cos_dat = 16'b1000101110001110;  
    10'd444     : cos_dat = 16'b1000101100111100;  
    10'd445     : cos_dat = 16'b1000101011101100;  
    10'd446     : cos_dat = 16'b1000101010011100;  
    10'd447     : cos_dat = 16'b1000101001001110;  
    10'd448     : cos_dat = 16'b1000101000000001;  
    10'd449     : cos_dat = 16'b1000100110110101;  
    10'd450     : cos_dat = 16'b1000100101101010;  
    10'd451     : cos_dat = 16'b1000100100100000;  
    10'd452     : cos_dat = 16'b1000100011011000;  
    10'd453     : cos_dat = 16'b1000100010010000;  
    10'd454     : cos_dat = 16'b1000100001001010;  
    10'd455     : cos_dat = 16'b1000100000000101;  
    10'd456     : cos_dat = 16'b1000011111000001;  
    10'd457     : cos_dat = 16'b1000011101111111;  
    10'd458     : cos_dat = 16'b1000011100111101;  
    10'd459     : cos_dat = 16'b1000011011111101;  
    10'd460     : cos_dat = 16'b1000011010111101;  
    10'd461     : cos_dat = 16'b1000011001111111;  
    10'd462     : cos_dat = 16'b1000011001000010;  
    10'd463     : cos_dat = 16'b1000011000000111;  
    10'd464     : cos_dat = 16'b1000010111001100;  
    10'd465     : cos_dat = 16'b1000010110010011;  
    10'd466     : cos_dat = 16'b1000010101011010;  
    10'd467     : cos_dat = 16'b1000010100100011;  
    10'd468     : cos_dat = 16'b1000010011101101;  
    10'd469     : cos_dat = 16'b1000010010111001;  
    10'd470     : cos_dat = 16'b1000010010000101;  
    10'd471     : cos_dat = 16'b1000010001010011;  
    10'd472     : cos_dat = 16'b1000010000100010;  
    10'd473     : cos_dat = 16'b1000001111110010;  
    10'd474     : cos_dat = 16'b1000001111000011;  
    10'd475     : cos_dat = 16'b1000001110010110;  
    10'd476     : cos_dat = 16'b1000001101101010;  
    10'd477     : cos_dat = 16'b1000001100111111;  
    10'd478     : cos_dat = 16'b1000001100010101;  
    10'd479     : cos_dat = 16'b1000001011101100;  
    10'd480     : cos_dat = 16'b1000001011000101;  
    10'd481     : cos_dat = 16'b1000001010011110;  
    10'd482     : cos_dat = 16'b1000001001111001;  
    10'd483     : cos_dat = 16'b1000001001010101;  
    10'd484     : cos_dat = 16'b1000001000110011;  
    10'd485     : cos_dat = 16'b1000001000010001;  
    10'd486     : cos_dat = 16'b1000000111110001;  
    10'd487     : cos_dat = 16'b1000000111010010;  
    10'd488     : cos_dat = 16'b1000000110110100;  
    10'd489     : cos_dat = 16'b1000000110011000;  
    10'd490     : cos_dat = 16'b1000000101111101;  
    10'd491     : cos_dat = 16'b1000000101100010;  
    10'd492     : cos_dat = 16'b1000000101001010;  
    10'd493     : cos_dat = 16'b1000000100110010;  
    10'd494     : cos_dat = 16'b1000000100011100;  
    10'd495     : cos_dat = 16'b1000000100000110;  
    10'd496     : cos_dat = 16'b1000000011110010;  
    10'd497     : cos_dat = 16'b1000000011100000;  
    10'd498     : cos_dat = 16'b1000000011001110;  
    10'd499     : cos_dat = 16'b1000000010111110;  
    10'd500     : cos_dat = 16'b1000000010101111;  
    10'd501     : cos_dat = 16'b1000000010100001;  
    10'd502     : cos_dat = 16'b1000000010010100;  
    10'd503     : cos_dat = 16'b1000000010001001;  
    10'd504     : cos_dat = 16'b1000000001111111;  
    10'd505     : cos_dat = 16'b1000000001110110;  
    10'd506     : cos_dat = 16'b1000000001101110;  
    10'd507     : cos_dat = 16'b1000000001100111;  
    10'd508     : cos_dat = 16'b1000000001100010;  
    10'd509     : cos_dat = 16'b1000000001011110;  
    10'd510     : cos_dat = 16'b1000000001011011;  
    10'd511     : cos_dat = 16'b1000000001011010;  
    10'd512     : cos_dat = 16'b1000000001011010;   
    10'd513     : cos_dat = 16'b1000000001011010;   
    10'd514     : cos_dat = 16'b1000000001011101;   
    10'd515     : cos_dat = 16'b1000000001100000;   
    10'd516     : cos_dat = 16'b1000000001100101;   
    10'd517     : cos_dat = 16'b1000000001101010;   
    10'd518     : cos_dat = 16'b1000000001110001;   
    10'd519     : cos_dat = 16'b1000000001111010;   
    10'd520     : cos_dat = 16'b1000000010000011;   
    10'd521     : cos_dat = 16'b1000000010001110;   
    10'd522     : cos_dat = 16'b1000000010011010;   
    10'd523     : cos_dat = 16'b1000000010100111;   
    10'd524     : cos_dat = 16'b1000000010110110;   
    10'd525     : cos_dat = 16'b1000000011000101;   
    10'd526     : cos_dat = 16'b1000000011010110;   
    10'd527     : cos_dat = 16'b1000000011101000;   
    10'd528     : cos_dat = 16'b1000000011111100;   
    10'd529     : cos_dat = 16'b1000000100010000;   
    10'd530     : cos_dat = 16'b1000000100100110;   
    10'd531     : cos_dat = 16'b1000000100111101;   
    10'd532     : cos_dat = 16'b1000000101010101;   
    10'd533     : cos_dat = 16'b1000000101101111;   
    10'd534     : cos_dat = 16'b1000000110001010;   
    10'd535     : cos_dat = 16'b1000000110100110;   
    10'd536     : cos_dat = 16'b1000000111000011;   
    10'd537     : cos_dat = 16'b1000000111100001;   
    10'd538     : cos_dat = 16'b1000001000000001;   
    10'd539     : cos_dat = 16'b1000001000100001;   
    10'd540     : cos_dat = 16'b1000001001000011;   
    10'd541     : cos_dat = 16'b1000001001100111;   
    10'd542     : cos_dat = 16'b1000001010001011;   
    10'd543     : cos_dat = 16'b1000001010110001;   
    10'd544     : cos_dat = 16'b1000001011010111;   
    10'd545     : cos_dat = 16'b1000001011111111;   
    10'd546     : cos_dat = 16'b1000001100101001;   
    10'd547     : cos_dat = 16'b1000001101010011;   
    10'd548     : cos_dat = 16'b1000001101111111;   
    10'd549     : cos_dat = 16'b1000001110101100;   
    10'd550     : cos_dat = 16'b1000001111011010;   
    10'd551     : cos_dat = 16'b1000010000001001;   
    10'd552     : cos_dat = 16'b1000010000111010;   
    10'd553     : cos_dat = 16'b1000010001101011;   
    10'd554     : cos_dat = 16'b1000010010011110;   
    10'd555     : cos_dat = 16'b1000010011010010;   
    10'd556     : cos_dat = 16'b1000010100000111;   
    10'd557     : cos_dat = 16'b1000010100111110;   
    10'd558     : cos_dat = 16'b1000010101110101;   
    10'd559     : cos_dat = 16'b1000010110101110;   
    10'd560     : cos_dat = 16'b1000010111101000;   
    10'd561     : cos_dat = 16'b1000011000100011;   
    10'd562     : cos_dat = 16'b1000011001011111;   
    10'd563     : cos_dat = 16'b1000011010011101;   
    10'd564     : cos_dat = 16'b1000011011011100;   
    10'd565     : cos_dat = 16'b1000011100011011;   
    10'd566     : cos_dat = 16'b1000011101011100;   
    10'd567     : cos_dat = 16'b1000011110011110;   
    10'd568     : cos_dat = 16'b1000011111100010;   
    10'd569     : cos_dat = 16'b1000100000100110;   
    10'd570     : cos_dat = 16'b1000100001101100;   
    10'd571     : cos_dat = 16'b1000100010110011;   
    10'd572     : cos_dat = 16'b1000100011111011;   
    10'd573     : cos_dat = 16'b1000100101000100;   
    10'd574     : cos_dat = 16'b1000100110001110;   
    10'd575     : cos_dat = 16'b1000100111011001;   
    10'd576     : cos_dat = 16'b1000101000100110;   
    10'd577     : cos_dat = 16'b1000101001110011;   
    10'd578     : cos_dat = 16'b1000101011000010;   
    10'd579     : cos_dat = 16'b1000101100010010;   
    10'd580     : cos_dat = 16'b1000101101100011;   
    10'd581     : cos_dat = 16'b1000101110110101;   
    10'd582     : cos_dat = 16'b1000110000001001;   
    10'd583     : cos_dat = 16'b1000110001011101;   
    10'd584     : cos_dat = 16'b1000110010110011;   
    10'd585     : cos_dat = 16'b1000110100001001;   
    10'd586     : cos_dat = 16'b1000110101100001;   
    10'd587     : cos_dat = 16'b1000110110111010;   
    10'd588     : cos_dat = 16'b1000111000010100;   
    10'd589     : cos_dat = 16'b1000111001101111;   
    10'd590     : cos_dat = 16'b1000111011001011;   
    10'd591     : cos_dat = 16'b1000111100101000;   
    10'd592     : cos_dat = 16'b1000111110000110;   
    10'd593     : cos_dat = 16'b1000111111100110;   
    10'd594     : cos_dat = 16'b1001000001000110;   
    10'd595     : cos_dat = 16'b1001000010101000;   
    10'd596     : cos_dat = 16'b1001000100001011;   
    10'd597     : cos_dat = 16'b1001000101101110;   
    10'd598     : cos_dat = 16'b1001000111010011;   
    10'd599     : cos_dat = 16'b1001001000111001;   
    10'd600     : cos_dat = 16'b1001001010100000;   
    10'd601     : cos_dat = 16'b1001001100001000;   
    10'd602     : cos_dat = 16'b1001001101110001;   
    10'd603     : cos_dat = 16'b1001001111011011;   
    10'd604     : cos_dat = 16'b1001010001000110;   
    10'd605     : cos_dat = 16'b1001010010110010;   
    10'd606     : cos_dat = 16'b1001010100011111;   
    10'd607     : cos_dat = 16'b1001010110001101;   
    10'd608     : cos_dat = 16'b1001010111111101;   
    10'd609     : cos_dat = 16'b1001011001101101;   
    10'd610     : cos_dat = 16'b1001011011011110;   
    10'd611     : cos_dat = 16'b1001011101010000;   
    10'd612     : cos_dat = 16'b1001011111000100;   
    10'd613     : cos_dat = 16'b1001100000111000;   
    10'd614     : cos_dat = 16'b1001100010101101;   
    10'd615     : cos_dat = 16'b1001100100100100;   
    10'd616     : cos_dat = 16'b1001100110011011;   
    10'd617     : cos_dat = 16'b1001101000010011;   
    10'd618     : cos_dat = 16'b1001101010001100;   
    10'd619     : cos_dat = 16'b1001101100000111;   
    10'd620     : cos_dat = 16'b1001101110000010;   
    10'd621     : cos_dat = 16'b1001101111111110;   
    10'd622     : cos_dat = 16'b1001110001111011;   
    10'd623     : cos_dat = 16'b1001110011111001;   
    10'd624     : cos_dat = 16'b1001110101111000;   
    10'd625     : cos_dat = 16'b1001110111111000;   
    10'd626     : cos_dat = 16'b1001111001111001;   
    10'd627     : cos_dat = 16'b1001111011111011;   
    10'd628     : cos_dat = 16'b1001111101111110;   
    10'd629     : cos_dat = 16'b1010000000000010;   
    10'd630     : cos_dat = 16'b1010000010000111;   
    10'd631     : cos_dat = 16'b1010000100001100;   
    10'd632     : cos_dat = 16'b1010000110010011;   
    10'd633     : cos_dat = 16'b1010001000011010;   
    10'd634     : cos_dat = 16'b1010001010100011;   
    10'd635     : cos_dat = 16'b1010001100101100;   
    10'd636     : cos_dat = 16'b1010001110110110;   
    10'd637     : cos_dat = 16'b1010010001000001;   
    10'd638     : cos_dat = 16'b1010010011001101;   
    10'd639     : cos_dat = 16'b1010010101011010;   
    10'd640     : cos_dat = 16'b1010010111100111;   
    10'd641     : cos_dat = 16'b1010011001110110;   
    10'd642     : cos_dat = 16'b1010011100000101;   
    10'd643     : cos_dat = 16'b1010011110010110;   
    10'd644     : cos_dat = 16'b1010100000100111;   
    10'd645     : cos_dat = 16'b1010100010111001;   
    10'd646     : cos_dat = 16'b1010100101001011;   
    10'd647     : cos_dat = 16'b1010100111011111;   
    10'd648     : cos_dat = 16'b1010101001110100;   
    10'd649     : cos_dat = 16'b1010101100001001;   
    10'd650     : cos_dat = 16'b1010101110011111;   
    10'd651     : cos_dat = 16'b1010110000110110;   
    10'd652     : cos_dat = 16'b1010110011001110;   
    10'd653     : cos_dat = 16'b1010110101100110;   
    10'd654     : cos_dat = 16'b1010111000000000;   
    10'd655     : cos_dat = 16'b1010111010011010;   
    10'd656     : cos_dat = 16'b1010111100110101;   
    10'd657     : cos_dat = 16'b1010111111010000;   
    10'd658     : cos_dat = 16'b1011000001101101;   
    10'd659     : cos_dat = 16'b1011000100001010;   
    10'd660     : cos_dat = 16'b1011000110101000;   
    10'd661     : cos_dat = 16'b1011001001000111;   
    10'd662     : cos_dat = 16'b1011001011100110;   
    10'd663     : cos_dat = 16'b1011001110000111;   
    10'd664     : cos_dat = 16'b1011010000101000;   
    10'd665     : cos_dat = 16'b1011010011001001;   
    10'd666     : cos_dat = 16'b1011010101101100;   
    10'd667     : cos_dat = 16'b1011011000001111;   
    10'd668     : cos_dat = 16'b1011011010110011;   
    10'd669     : cos_dat = 16'b1011011101010111;   
    10'd670     : cos_dat = 16'b1011011111111101;   
    10'd671     : cos_dat = 16'b1011100010100011;   
    10'd672     : cos_dat = 16'b1011100101001001;   
    10'd673     : cos_dat = 16'b1011100111110001;   
    10'd674     : cos_dat = 16'b1011101010011001;   
    10'd675     : cos_dat = 16'b1011101101000001;   
    10'd676     : cos_dat = 16'b1011101111101011;   
    10'd677     : cos_dat = 16'b1011110010010101;   
    10'd678     : cos_dat = 16'b1011110100111111;   
    10'd679     : cos_dat = 16'b1011110111101011;   
    10'd680     : cos_dat = 16'b1011111010010111;   
    10'd681     : cos_dat = 16'b1011111101000011;   
    10'd682     : cos_dat = 16'b1011111111110000;   
    10'd683     : cos_dat = 16'b1100000010011110;   
    10'd684     : cos_dat = 16'b1100000101001101;   
    10'd685     : cos_dat = 16'b1100000111111100;   
    10'd686     : cos_dat = 16'b1100001010101011;   
    10'd687     : cos_dat = 16'b1100001101011100;   
    10'd688     : cos_dat = 16'b1100010000001100;   
    10'd689     : cos_dat = 16'b1100010010111110;   
    10'd690     : cos_dat = 16'b1100010101110000;   
    10'd691     : cos_dat = 16'b1100011000100010;   
    10'd692     : cos_dat = 16'b1100011011010101;   
    10'd693     : cos_dat = 16'b1100011110001001;   
    10'd694     : cos_dat = 16'b1100100000111101;   
    10'd695     : cos_dat = 16'b1100100011110010;   
    10'd696     : cos_dat = 16'b1100100110100111;   
    10'd697     : cos_dat = 16'b1100101001011101;   
    10'd698     : cos_dat = 16'b1100101100010011;   
    10'd699     : cos_dat = 16'b1100101111001010;   
    10'd700     : cos_dat = 16'b1100110010000001;   
    10'd701     : cos_dat = 16'b1100110100111001;   
    10'd702     : cos_dat = 16'b1100110111110001;   
    10'd703     : cos_dat = 16'b1100111010101010;   
    10'd704     : cos_dat = 16'b1100111101100011;   
    10'd705     : cos_dat = 16'b1101000000011101;   
    10'd706     : cos_dat = 16'b1101000011010111;   
    10'd707     : cos_dat = 16'b1101000110010010;   
    10'd708     : cos_dat = 16'b1101001001001101;   
    10'd709     : cos_dat = 16'b1101001100001001;   
    10'd710     : cos_dat = 16'b1101001111000101;   
    10'd711     : cos_dat = 16'b1101010010000001;   
    10'd712     : cos_dat = 16'b1101010100111110;   
    10'd713     : cos_dat = 16'b1101010111111011;   
    10'd714     : cos_dat = 16'b1101011010111001;   
    10'd715     : cos_dat = 16'b1101011101110111;   
    10'd716     : cos_dat = 16'b1101100000110101;   
    10'd717     : cos_dat = 16'b1101100011110100;   
    10'd718     : cos_dat = 16'b1101100110110011;   
    10'd719     : cos_dat = 16'b1101101001110011;   
    10'd720     : cos_dat = 16'b1101101100110011;   
    10'd721     : cos_dat = 16'b1101101111110011;   
    10'd722     : cos_dat = 16'b1101110010110011;   
    10'd723     : cos_dat = 16'b1101110101110100;   
    10'd724     : cos_dat = 16'b1101111000110110;   
    10'd725     : cos_dat = 16'b1101111011110111;   
    10'd726     : cos_dat = 16'b1101111110111001;   
    10'd727     : cos_dat = 16'b1110000001111011;   
    10'd728     : cos_dat = 16'b1110000100111110;   
    10'd729     : cos_dat = 16'b1110001000000001;   
    10'd730     : cos_dat = 16'b1110001011000100;   
    10'd731     : cos_dat = 16'b1110001110000111;   
    10'd732     : cos_dat = 16'b1110010001001011;   
    10'd733     : cos_dat = 16'b1110010100001111;   
    10'd734     : cos_dat = 16'b1110010111010011;   
    10'd735     : cos_dat = 16'b1110011010011000;   
    10'd736     : cos_dat = 16'b1110011101011100;   
    10'd737     : cos_dat = 16'b1110100000100001;   
    10'd738     : cos_dat = 16'b1110100011100111;   
    10'd739     : cos_dat = 16'b1110100110101100;   
    10'd740     : cos_dat = 16'b1110101001110010;   
    10'd741     : cos_dat = 16'b1110101100110111;   
    10'd742     : cos_dat = 16'b1110101111111101;   
    10'd743     : cos_dat = 16'b1110110011000100;   
    10'd744     : cos_dat = 16'b1110110110001010;   
    10'd745     : cos_dat = 16'b1110111001010001;   
    10'd746     : cos_dat = 16'b1110111100010111;   
    10'd747     : cos_dat = 16'b1110111111011110;   
    10'd748     : cos_dat = 16'b1111000010100101;   
    10'd749     : cos_dat = 16'b1111000101101101;   
    10'd750     : cos_dat = 16'b1111001000110100;   
    10'd751     : cos_dat = 16'b1111001011111011;   
    10'd752     : cos_dat = 16'b1111001111000011;   
    10'd753     : cos_dat = 16'b1111010010001011;   
    10'd754     : cos_dat = 16'b1111010101010011;   
    10'd755     : cos_dat = 16'b1111011000011011;   
    10'd756     : cos_dat = 16'b1111011011100011;   
    10'd757     : cos_dat = 16'b1111011110101011;   
    10'd758     : cos_dat = 16'b1111100001110011;   
    10'd759     : cos_dat = 16'b1111100100111011;   
    10'd760     : cos_dat = 16'b1111101000000100;   
    10'd761     : cos_dat = 16'b1111101011001100;   
    10'd762     : cos_dat = 16'b1111101110010100;   
    10'd763     : cos_dat = 16'b1111110001011101;   
    10'd764     : cos_dat = 16'b1111110100100110;   
    10'd765     : cos_dat = 16'b1111110111101110;   
    10'd766     : cos_dat = 16'b1111111010110111;   
    10'd767     : cos_dat = 16'b1111111101111111;   
    10'd768     : cos_dat = 16'b0000000001001000;   
    10'd769     : cos_dat = 16'b0000000100010000;   
    10'd770     : cos_dat = 16'b0000000111011001;   
    10'd771     : cos_dat = 16'b0000001010100010;   
    10'd772     : cos_dat = 16'b0000001101101010;   
    10'd773     : cos_dat = 16'b0000010000110011;   
    10'd774     : cos_dat = 16'b0000010011111011;   
    10'd775     : cos_dat = 16'b0000010111000100;   
    10'd776     : cos_dat = 16'b0000011010001100;   
    10'd777     : cos_dat = 16'b0000011101010100;   
    10'd778     : cos_dat = 16'b0000100000011101;   
    10'd779     : cos_dat = 16'b0000100011100101;   
    10'd780     : cos_dat = 16'b0000100110101101;   
    10'd781     : cos_dat = 16'b0000101001110101;   
    10'd782     : cos_dat = 16'b0000101100111101;   
    10'd783     : cos_dat = 16'b0000110000000100;   
    10'd784     : cos_dat = 16'b0000110011001100;   
    10'd785     : cos_dat = 16'b0000110110010100;   
    10'd786     : cos_dat = 16'b0000111001011011;   
    10'd787     : cos_dat = 16'b0000111100100010;   
    10'd788     : cos_dat = 16'b0000111111101001;   
    10'd789     : cos_dat = 16'b0001000010110000;   
    10'd790     : cos_dat = 16'b0001000101110111;   
    10'd791     : cos_dat = 16'b0001001000111110;   
    10'd792     : cos_dat = 16'b0001001100000100;   
    10'd793     : cos_dat = 16'b0001001111001010;   
    10'd794     : cos_dat = 16'b0001010010010001;   
    10'd795     : cos_dat = 16'b0001010101010110;   
    10'd796     : cos_dat = 16'b0001011000011100;   
    10'd797     : cos_dat = 16'b0001011011100010;   
    10'd798     : cos_dat = 16'b0001011110100111;   
    10'd799     : cos_dat = 16'b0001100001101100;   
    10'd800     : cos_dat = 16'b0001100100110001;   
    10'd801     : cos_dat = 16'b0001100111110101;   
    10'd802     : cos_dat = 16'b0001101010111001;   
    10'd803     : cos_dat = 16'b0001101101111101;   
    10'd804     : cos_dat = 16'b0001110001000001;   
    10'd805     : cos_dat = 16'b0001110100000101;   
    10'd806     : cos_dat = 16'b0001110111001000;   
    10'd807     : cos_dat = 16'b0001111010001011;   
    10'd808     : cos_dat = 16'b0001111101001101;   
    10'd809     : cos_dat = 16'b0010000000010000;   
    10'd810     : cos_dat = 16'b0010000011010010;   
    10'd811     : cos_dat = 16'b0010000110010100;   
    10'd812     : cos_dat = 16'b0010001001010101;   
    10'd813     : cos_dat = 16'b0010001100010110;   
    10'd814     : cos_dat = 16'b0010001111010111;   
    10'd815     : cos_dat = 16'b0010010010010111;   
    10'd816     : cos_dat = 16'b0010010101010111;   
    10'd817     : cos_dat = 16'b0010011000010111;   
    10'd818     : cos_dat = 16'b0010011011010110;   
    10'd819     : cos_dat = 16'b0010011110010101;   
    10'd820     : cos_dat = 16'b0010100001010011;   
    10'd821     : cos_dat = 16'b0010100100010001;   
    10'd822     : cos_dat = 16'b0010100111001111;   
    10'd823     : cos_dat = 16'b0010101010001101;   
    10'd824     : cos_dat = 16'b0010101101001001;   
    10'd825     : cos_dat = 16'b0010110000000110;   
    10'd826     : cos_dat = 16'b0010110011000010;   
    10'd827     : cos_dat = 16'b0010110101111110;   
    10'd828     : cos_dat = 16'b0010111000111001;   
    10'd829     : cos_dat = 16'b0010111011110100;   
    10'd830     : cos_dat = 16'b0010111110101110;   
    10'd831     : cos_dat = 16'b0011000001101000;   
    10'd832     : cos_dat = 16'b0011000100100001;   
    10'd833     : cos_dat = 16'b0011000111011010;   
    10'd834     : cos_dat = 16'b0011001010010011;   
    10'd835     : cos_dat = 16'b0011001101001011;   
    10'd836     : cos_dat = 16'b0011010000000010;   
    10'd837     : cos_dat = 16'b0011010010111001;   
    10'd838     : cos_dat = 16'b0011010101101111;   
    10'd839     : cos_dat = 16'b0011011000100101;   
    10'd840     : cos_dat = 16'b0011011011011011;   
    10'd841     : cos_dat = 16'b0011011110010000;   
    10'd842     : cos_dat = 16'b0011100001000100;   
    10'd843     : cos_dat = 16'b0011100011111000;   
    10'd844     : cos_dat = 16'b0011100110101011;   
    10'd845     : cos_dat = 16'b0011101001011110;   
    10'd846     : cos_dat = 16'b0011101100010000;   
    10'd847     : cos_dat = 16'b0011101111000001;   
    10'd848     : cos_dat = 16'b0011110001110010;   
    10'd849     : cos_dat = 16'b0011110100100011;   
    10'd850     : cos_dat = 16'b0011110111010010;   
    10'd851     : cos_dat = 16'b0011111010000010;   
    10'd852     : cos_dat = 16'b0011111100110000;   
    10'd853     : cos_dat = 16'b0011111111011110;   
    10'd854     : cos_dat = 16'b0100000010001100;   
    10'd855     : cos_dat = 16'b0100000100111000;   
    10'd856     : cos_dat = 16'b0100000111100100;   
    10'd857     : cos_dat = 16'b0100001010010000;   
    10'd858     : cos_dat = 16'b0100001100111011;   
    10'd859     : cos_dat = 16'b0100001111100101;   
    10'd860     : cos_dat = 16'b0100010010001111;   
    10'd861     : cos_dat = 16'b0100010100110111;   
    10'd862     : cos_dat = 16'b0100010111100000;   
    10'd863     : cos_dat = 16'b0100011010000111;   
    10'd864     : cos_dat = 16'b0100011100101110;   
    10'd865     : cos_dat = 16'b0100011111010100;   
    10'd866     : cos_dat = 16'b0100100001111010;   
    10'd867     : cos_dat = 16'b0100100100011111;   
    10'd868     : cos_dat = 16'b0100100111000011;   
    10'd869     : cos_dat = 16'b0100101001100110;   
    10'd870     : cos_dat = 16'b0100101100001001;   
    10'd871     : cos_dat = 16'b0100101110101011;   
    10'd872     : cos_dat = 16'b0100110001001100;   
    10'd873     : cos_dat = 16'b0100110011101100;   
    10'd874     : cos_dat = 16'b0100110110001100;   
    10'd875     : cos_dat = 16'b0100111000101011;   
    10'd876     : cos_dat = 16'b0100111011001001;   
    10'd877     : cos_dat = 16'b0100111101100111;   
    10'd878     : cos_dat = 16'b0101000000000011;   
    10'd879     : cos_dat = 16'b0101000010011111;   
    10'd880     : cos_dat = 16'b0101000100111010;   
    10'd881     : cos_dat = 16'b0101000111010101;   
    10'd882     : cos_dat = 16'b0101001001101110;   
    10'd883     : cos_dat = 16'b0101001100000111;   
    10'd884     : cos_dat = 16'b0101001110011111;   
    10'd885     : cos_dat = 16'b0101010000110110;   
    10'd886     : cos_dat = 16'b0101010011001100;   
    10'd887     : cos_dat = 16'b0101010101100010;   
    10'd888     : cos_dat = 16'b0101010111110111;   
    10'd889     : cos_dat = 16'b0101011010001011;   
    10'd890     : cos_dat = 16'b0101011100011110;   
    10'd891     : cos_dat = 16'b0101011110110000;   
    10'd892     : cos_dat = 16'b0101100001000001;   
    10'd893     : cos_dat = 16'b0101100011010010;   
    10'd894     : cos_dat = 16'b0101100101100001;   
    10'd895     : cos_dat = 16'b0101100111110000;   
    10'd896     : cos_dat = 16'b0101101001111110;   
    10'd897     : cos_dat = 16'b0101101100001011;   
    10'd898     : cos_dat = 16'b0101101110010111;   
    10'd899     : cos_dat = 16'b0101110000100010;   
    10'd900     : cos_dat = 16'b0101110010101101;   
    10'd901     : cos_dat = 16'b0101110100110110;   
    10'd902     : cos_dat = 16'b0101110110111111;   
    10'd903     : cos_dat = 16'b0101111001000111;   
    10'd904     : cos_dat = 16'b0101111011001101;   
    10'd905     : cos_dat = 16'b0101111101010011;   
    10'd906     : cos_dat = 16'b0101111111011000;   
    10'd907     : cos_dat = 16'b0110000001011100;   
    10'd908     : cos_dat = 16'b0110000011011111;   
    10'd909     : cos_dat = 16'b0110000101100010;   
    10'd910     : cos_dat = 16'b0110000111100011;   
    10'd911     : cos_dat = 16'b0110001001100011;   
    10'd912     : cos_dat = 16'b0110001011100010;   
    10'd913     : cos_dat = 16'b0110001101100001;   
    10'd914     : cos_dat = 16'b0110001111011110;   
    10'd915     : cos_dat = 16'b0110010001011011;   
    10'd916     : cos_dat = 16'b0110010011010110;   
    10'd917     : cos_dat = 16'b0110010101010001;   
    10'd918     : cos_dat = 16'b0110010111001010;   
    10'd919     : cos_dat = 16'b0110011001000011;   
    10'd920     : cos_dat = 16'b0110011010111010;   
    10'd921     : cos_dat = 16'b0110011100110001;   
    10'd922     : cos_dat = 16'b0110011110100110;   
    10'd923     : cos_dat = 16'b0110100000011011;   
    10'd924     : cos_dat = 16'b0110100010001111;   
    10'd925     : cos_dat = 16'b0110100100000001;   
    10'd926     : cos_dat = 16'b0110100101110011;   
    10'd927     : cos_dat = 16'b0110100111100011;   
    10'd928     : cos_dat = 16'b0110101001010011;   
    10'd929     : cos_dat = 16'b0110101011000001;   
    10'd930     : cos_dat = 16'b0110101100101111;   
    10'd931     : cos_dat = 16'b0110101110011011;   
    10'd932     : cos_dat = 16'b0110110000000111;   
    10'd933     : cos_dat = 16'b0110110001110001;   
    10'd934     : cos_dat = 16'b0110110011011010;   
    10'd935     : cos_dat = 16'b0110110101000010;   
    10'd936     : cos_dat = 16'b0110110110101010;   
    10'd937     : cos_dat = 16'b0110111000010000;   
    10'd938     : cos_dat = 16'b0110111001110101;   
    10'd939     : cos_dat = 16'b0110111011011001;   
    10'd940     : cos_dat = 16'b0110111100111100;   
    10'd941     : cos_dat = 16'b0110111110011110;   
    10'd942     : cos_dat = 16'b0110111111111110;   
    10'd943     : cos_dat = 16'b0111000001011110;   
    10'd944     : cos_dat = 16'b0111000010111101;   
    10'd945     : cos_dat = 16'b0111000100011010;   
    10'd946     : cos_dat = 16'b0111000101110111;   
    10'd947     : cos_dat = 16'b0111000111010010;   
    10'd948     : cos_dat = 16'b0111001000101100;   
    10'd949     : cos_dat = 16'b0111001010000110;   
    10'd950     : cos_dat = 16'b0111001011011110;   
    10'd951     : cos_dat = 16'b0111001100110100;   
    10'd952     : cos_dat = 16'b0111001110001010;   
    10'd953     : cos_dat = 16'b0111001111011111;   
    10'd954     : cos_dat = 16'b0111010000110011;   
    10'd955     : cos_dat = 16'b0111010010000101;   
    10'd956     : cos_dat = 16'b0111010011010110;   
    10'd957     : cos_dat = 16'b0111010100100111;   
    10'd958     : cos_dat = 16'b0111010101110110;   
    10'd959     : cos_dat = 16'b0111010111000100;   
    10'd960     : cos_dat = 16'b0111011000010001;   
    10'd961     : cos_dat = 16'b0111011001011100;   
    10'd962     : cos_dat = 16'b0111011010100111;   
    10'd963     : cos_dat = 16'b0111011011110000;   
    10'd964     : cos_dat = 16'b0111011100111000;   
    10'd965     : cos_dat = 16'b0111011110000000;   
    10'd966     : cos_dat = 16'b0111011111000101;   
    10'd967     : cos_dat = 16'b0111100000001010;   
    10'd968     : cos_dat = 16'b0111100001001110;   
    10'd969     : cos_dat = 16'b0111100010010000;   
    10'd970     : cos_dat = 16'b0111100011010010;   
    10'd971     : cos_dat = 16'b0111100100010010;   
    10'd972     : cos_dat = 16'b0111100101010001;   
    10'd973     : cos_dat = 16'b0111100110001111;   
    10'd974     : cos_dat = 16'b0111100111001011;   
    10'd975     : cos_dat = 16'b0111101000000111;   
    10'd976     : cos_dat = 16'b0111101001000001;   
    10'd977     : cos_dat = 16'b0111101001111010;   
    10'd978     : cos_dat = 16'b0111101010110010;   
    10'd979     : cos_dat = 16'b0111101011101001;   
    10'd980     : cos_dat = 16'b0111101100011110;   
    10'd981     : cos_dat = 16'b0111101101010011;   
    10'd982     : cos_dat = 16'b0111101110000110;   
    10'd983     : cos_dat = 16'b0111101110111000;   
    10'd984     : cos_dat = 16'b0111101111101001;   
    10'd985     : cos_dat = 16'b0111110000011000;   
    10'd986     : cos_dat = 16'b0111110001000111;   
    10'd987     : cos_dat = 16'b0111110001110100;   
    10'd988     : cos_dat = 16'b0111110010100000;   
    10'd989     : cos_dat = 16'b0111110011001011;   
    10'd990     : cos_dat = 16'b0111110011110100;   
    10'd991     : cos_dat = 16'b0111110100011101;   
    10'd992     : cos_dat = 16'b0111110101000100;   
    10'd993     : cos_dat = 16'b0111110101101010;   
    10'd994     : cos_dat = 16'b0111110110001110;   
    10'd995     : cos_dat = 16'b0111110110110010;   
    10'd996     : cos_dat = 16'b0111110111010100;   
    10'd997     : cos_dat = 16'b0111110111110101;   
    10'd998     : cos_dat = 16'b0111111000010101;   
    10'd999     : cos_dat = 16'b0111111000110100;   
    10'd1000    : cos_dat = 16'b0111111001010010;   
    10'd1001    : cos_dat = 16'b0111111001101110;   
    10'd1002    : cos_dat = 16'b0111111010001001;   
    10'd1003    : cos_dat = 16'b0111111010100011;   
    10'd1004    : cos_dat = 16'b0111111010111011;   
    10'd1005    : cos_dat = 16'b0111111011010011;   
    10'd1006    : cos_dat = 16'b0111111011101001;   
    10'd1007    : cos_dat = 16'b0111111011111110;   
    10'd1008    : cos_dat = 16'b0111111100010001;   
    10'd1009    : cos_dat = 16'b0111111100100100;   
    10'd1010    : cos_dat = 16'b0111111100110101;   
    10'd1011    : cos_dat = 16'b0111111101000101;   
    10'd1012    : cos_dat = 16'b0111111101010100;   
    10'd1013    : cos_dat = 16'b0111111101100001;   
    10'd1014    : cos_dat = 16'b0111111101101110;   
    10'd1015    : cos_dat = 16'b0111111101111001;   
    10'd1016    : cos_dat = 16'b0111111110000011;   
    10'd1017    : cos_dat = 16'b0111111110001011;   
    10'd1018    : cos_dat = 16'b0111111110010011;   
    10'd1019    : cos_dat = 16'b0111111110011001;   
    10'd1020    : cos_dat = 16'b0111111110011110;   
    10'd1021    : cos_dat = 16'b0111111110100010;   
    10'd1022    : cos_dat = 16'b0111111110100100;   
    10'd1023    : cos_dat = 16'b0111111110100101;   
    default     : cos_dat = 16'b0000000000000000;  
    endcase
end



//*******************************************************************************
//
// END of Module
//
//*******************************************************************************
endmodule
