
class ral_reg_HOST_ID extends uvm_reg;



endclass




