
`timescale 1ns / 1ps

//--------------------------
// rtl
//--------------------------
`include "../rtl/router.sv"

//--------------------------
// interface
//--------------------------
`include "router_io.sv"



//----------------------------------------------------------//
//
// testbench
//
//----------------------------------------------------------//
module top;








endmodule
//----------------------------------------------------------//
//
// End of Module
//
//----------------------------------------------------------//

