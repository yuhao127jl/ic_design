//*******************************************************************************
// Project      : 
// Module       : rs_lat.v
// Description  :
// Designer     :
// Version      : 
//********************************************************************************

module rs_lat(
input  wire     rn,
input  wire     sn,
output wire     q,
output wire     qn
);


NAND2HD2X nd0(.A(rn), .B(q),  .Z(qn));
NAND2HD2X nd1(.A(rn), .B(qn), .Z(q));



//********************************************************************************
//
// END of Module
//
//********************************************************************************
endmodule
