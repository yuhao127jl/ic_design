//*******************************************************************************
// Project		: 
// Module		: sin_tbl.v
// Description	: 
// Designer		: 
// Version		: 
//*******************************************************************************

module sin_tbl(
    input wire[9:0]      addr,
    output reg[15:0]     sin_dat
);

//**********************************************************
//
// always
//
//**********************************************************
always @(*)
begin
    case(addr)
    10'd0       : sin_dat = 16'b0000000000000000 ;  
    10'd1       : sin_dat = 16'b0000000011001000 ;  
    10'd2       : sin_dat = 16'b0000000110010001 ;  
    10'd3       : sin_dat = 16'b0000001001011001 ;  
    10'd4       : sin_dat = 16'b0000001100100010 ;  
    10'd5       : sin_dat = 16'b0000001111101010 ;  
    10'd6       : sin_dat = 16'b0000010010110011 ;  
    10'd7       : sin_dat = 16'b0000010101111011 ;  
    10'd8       : sin_dat = 16'b0000011001000100 ;  
    10'd9       : sin_dat = 16'b0000011100001100 ;  
    10'd10      : sin_dat = 16'b0000011111010100 ;  
    10'd11      : sin_dat = 16'b0000100010011100 ;  
    10'd12      : sin_dat = 16'b0000100101100101 ;  
    10'd13      : sin_dat = 16'b0000101000101101 ;  
    10'd14      : sin_dat = 16'b0000101011110100 ;  
    10'd15      : sin_dat = 16'b0000101110111100 ;  
    10'd16      : sin_dat = 16'b0000110010000100 ;  
    10'd17      : sin_dat = 16'b0000110101001100 ;  
    10'd18      : sin_dat = 16'b0000111000010011 ;  
    10'd19      : sin_dat = 16'b0000111011011010 ;  
    10'd20      : sin_dat = 16'b0000111110100010 ;  
    10'd21      : sin_dat = 16'b0001000001101001 ;  
    10'd22      : sin_dat = 16'b0001000100101111 ;  
    10'd23      : sin_dat = 16'b0001000111110110 ;  
    10'd24      : sin_dat = 16'b0001001010111101 ;  
    10'd25      : sin_dat = 16'b0001001110000011 ;  
    10'd26      : sin_dat = 16'b0001010001001001 ;  
    10'd27      : sin_dat = 16'b0001010100001111 ;  
    10'd28      : sin_dat = 16'b0001010111010101 ;  
    10'd29      : sin_dat = 16'b0001011010011010 ;  
    10'd30      : sin_dat = 16'b0001011101100000 ;  
    10'd31      : sin_dat = 16'b0001100000100101 ;  
    10'd32      : sin_dat = 16'b0001100011101010 ;  
    10'd33      : sin_dat = 16'b0001100110101110 ;  
    10'd34      : sin_dat = 16'b0001101001110011 ;  
    10'd35      : sin_dat = 16'b0001101100110111 ;  
    10'd36      : sin_dat = 16'b0001101111111011 ;  
    10'd37      : sin_dat = 16'b0001110010111110 ;  
    10'd38      : sin_dat = 16'b0001110110000010 ;  
    10'd39      : sin_dat = 16'b0001111001000101 ;  
    10'd40      : sin_dat = 16'b0001111100000111 ;  
    10'd41      : sin_dat = 16'b0001111111001010 ;  
    10'd42      : sin_dat = 16'b0010000010001100 ;  
    10'd43      : sin_dat = 16'b0010000101001110 ;  
    10'd44      : sin_dat = 16'b0010001000001111 ;  
    10'd45      : sin_dat = 16'b0010001011010000 ;  
    10'd46      : sin_dat = 16'b0010001110010001 ;  
    10'd47      : sin_dat = 16'b0010010001010010 ;  
    10'd48      : sin_dat = 16'b0010010100010010 ;  
    10'd49      : sin_dat = 16'b0010010111010010 ;  
    10'd50      : sin_dat = 16'b0010011010010001 ;  
    10'd51      : sin_dat = 16'b0010011101010000 ;  
    10'd52      : sin_dat = 16'b0010100000001111 ;  
    10'd53      : sin_dat = 16'b0010100011001101 ;  
    10'd54      : sin_dat = 16'b0010100110001011 ;  
    10'd55      : sin_dat = 16'b0010101001001000 ;  
    10'd56      : sin_dat = 16'b0010101100000101 ;  
    10'd57      : sin_dat = 16'b0010101111000010 ;  
    10'd58      : sin_dat = 16'b0010110001111110 ;  
    10'd59      : sin_dat = 16'b0010110100111010 ;  
    10'd60      : sin_dat = 16'b0010110111110101 ;  
    10'd61      : sin_dat = 16'b0010111010110000 ;  
    10'd62      : sin_dat = 16'b0010111101101011 ;  
    10'd63      : sin_dat = 16'b0011000000100101 ;  
    10'd64      : sin_dat = 16'b0011000011011110 ;  
    10'd65      : sin_dat = 16'b0011000110010111 ;  
    10'd66      : sin_dat = 16'b0011001001010000 ;  
    10'd67      : sin_dat = 16'b0011001100001000 ;  
    10'd68      : sin_dat = 16'b0011001111000000 ;  
    10'd69      : sin_dat = 16'b0011010001110111 ;  
    10'd70      : sin_dat = 16'b0011010100101110 ;  
    10'd71      : sin_dat = 16'b0011010111100100 ;  
    10'd72      : sin_dat = 16'b0011011010011001 ;  
    10'd73      : sin_dat = 16'b0011011101001110 ;  
    10'd74      : sin_dat = 16'b0011100000000011 ;  
    10'd75      : sin_dat = 16'b0011100010110111 ;  
    10'd76      : sin_dat = 16'b0011100101101010 ;  
    10'd77      : sin_dat = 16'b0011101000011101 ;  
    10'd78      : sin_dat = 16'b0011101011010000 ;  
    10'd79      : sin_dat = 16'b0011101110000001 ;  
    10'd80      : sin_dat = 16'b0011110000110010 ;  
    10'd81      : sin_dat = 16'b0011110011100011 ;  
    10'd82      : sin_dat = 16'b0011110110010011 ;  
    10'd83      : sin_dat = 16'b0011111001000010 ;  
    10'd84      : sin_dat = 16'b0011111011110001 ;  
    10'd85      : sin_dat = 16'b0011111110100000 ;  
    10'd86      : sin_dat = 16'b0100000001001101 ;  
    10'd87      : sin_dat = 16'b0100000011111010 ;  
    10'd88      : sin_dat = 16'b0100000110100110 ;  
    10'd89      : sin_dat = 16'b0100001001010010 ;  
    10'd90      : sin_dat = 16'b0100001011111101 ;  
    10'd91      : sin_dat = 16'b0100001110101000 ;  
    10'd92      : sin_dat = 16'b0100010001010001 ;  
    10'd93      : sin_dat = 16'b0100010011111011 ;  
    10'd94      : sin_dat = 16'b0100010110100011 ;  
    10'd95      : sin_dat = 16'b0100011001001011 ;  
    10'd96      : sin_dat = 16'b0100011011110010 ;  
    10'd97      : sin_dat = 16'b0100011110011000 ;  
    10'd98      : sin_dat = 16'b0100100000111110 ;  
    10'd99      : sin_dat = 16'b0100100011100011 ;  
    10'd100     : sin_dat = 16'b0100100110000111 ;  
    10'd101     : sin_dat = 16'b0100101000101011 ;  
    10'd102     : sin_dat = 16'b0100101011001110 ;  
    10'd103     : sin_dat = 16'b0100101101110000 ;  
    10'd104     : sin_dat = 16'b0100110000010010 ;  
    10'd105     : sin_dat = 16'b0100110010110010 ;  
    10'd106     : sin_dat = 16'b0100110101010010 ;  
    10'd107     : sin_dat = 16'b0100110111110010 ;  
    10'd108     : sin_dat = 16'b0100111010010000 ;  
    10'd109     : sin_dat = 16'b0100111100101110 ;  
    10'd110     : sin_dat = 16'b0100111111001011 ;  
    10'd111     : sin_dat = 16'b0101000001100111 ;  
    10'd112     : sin_dat = 16'b0101000100000010 ;  
    10'd113     : sin_dat = 16'b0101000110011101 ;  
    10'd114     : sin_dat = 16'b0101001000110111 ;  
    10'd115     : sin_dat = 16'b0101001011010000 ;  
    10'd116     : sin_dat = 16'b0101001101101000 ;  
    10'd117     : sin_dat = 16'b0101010000000000 ;  
    10'd118     : sin_dat = 16'b0101010010010110 ;  
    10'd119     : sin_dat = 16'b0101010100101100 ;  
    10'd120     : sin_dat = 16'b0101010111000001 ;  
    10'd121     : sin_dat = 16'b0101011001010101 ;  
    10'd122     : sin_dat = 16'b0101011011101001 ;  
    10'd123     : sin_dat = 16'b0101011101111011 ;  
    10'd124     : sin_dat = 16'b0101100000001101 ;  
    10'd125     : sin_dat = 16'b0101100010011110 ;  
    10'd126     : sin_dat = 16'b0101100100101110 ;  
    10'd127     : sin_dat = 16'b0101100110111101 ;  
    10'd128     : sin_dat = 16'b0101101001001011 ;  
    10'd129     : sin_dat = 16'b0101101011011000 ;  
    10'd130     : sin_dat = 16'b0101101101100101 ;  
    10'd131     : sin_dat = 16'b0101101111110000 ;  
    10'd132     : sin_dat = 16'b0101110001111011 ;  
    10'd133     : sin_dat = 16'b0101110100000101 ;  
    10'd134     : sin_dat = 16'b0101110110001110 ;  
    10'd135     : sin_dat = 16'b0101111000010110 ;  
    10'd136     : sin_dat = 16'b0101111010011101 ;  
    10'd137     : sin_dat = 16'b0101111100100011 ;  
    10'd138     : sin_dat = 16'b0101111110101000 ;  
    10'd139     : sin_dat = 16'b0110000000101101 ;  
    10'd140     : sin_dat = 16'b0110000010110000 ;  
    10'd141     : sin_dat = 16'b0110000100110011 ;  
    10'd142     : sin_dat = 16'b0110000110110100 ;  
    10'd143     : sin_dat = 16'b0110001000110101 ;  
    10'd144     : sin_dat = 16'b0110001010110101 ;  
    10'd145     : sin_dat = 16'b0110001100110011 ;  
    10'd146     : sin_dat = 16'b0110001110110001 ;  
    10'd147     : sin_dat = 16'b0110010000101110 ;  
    10'd148     : sin_dat = 16'b0110010010101010 ;  
    10'd149     : sin_dat = 16'b0110010100100101 ;  
    10'd150     : sin_dat = 16'b0110010110011110 ;  
    10'd151     : sin_dat = 16'b0110011000010111 ;  
    10'd152     : sin_dat = 16'b0110011010001111 ;  
    10'd153     : sin_dat = 16'b0110011100000110 ;  
    10'd154     : sin_dat = 16'b0110011101111100 ;  
    10'd155     : sin_dat = 16'b0110011111110001 ;  
    10'd156     : sin_dat = 16'b0110100001100101 ;  
    10'd157     : sin_dat = 16'b0110100011011000 ;  
    10'd158     : sin_dat = 16'b0110100101001010 ;  
    10'd159     : sin_dat = 16'b0110100110111011 ;  
    10'd160     : sin_dat = 16'b0110101000101011 ;  
    10'd161     : sin_dat = 16'b0110101010011001 ;  
    10'd162     : sin_dat = 16'b0110101100000111 ;  
    10'd163     : sin_dat = 16'b0110101101110100 ;  
    10'd164     : sin_dat = 16'b0110101111100000 ;  
    10'd165     : sin_dat = 16'b0110110001001011 ;  
    10'd166     : sin_dat = 16'b0110110010110100 ;  
    10'd167     : sin_dat = 16'b0110110100011101 ;  
    10'd168     : sin_dat = 16'b0110110110000100 ;  
    10'd169     : sin_dat = 16'b0110110111101011 ;  
    10'd170     : sin_dat = 16'b0110111001010000 ;  
    10'd171     : sin_dat = 16'b0110111010110101 ;  
    10'd172     : sin_dat = 16'b0110111100011000 ;  
    10'd173     : sin_dat = 16'b0110111101111010 ;  
    10'd174     : sin_dat = 16'b0110111111011100 ;  
    10'd175     : sin_dat = 16'b0111000000111100 ;  
    10'd176     : sin_dat = 16'b0111000010011011 ;  
    10'd177     : sin_dat = 16'b0111000011111001 ;  
    10'd178     : sin_dat = 16'b0111000101010110 ;  
    10'd179     : sin_dat = 16'b0111000110110001 ;  
    10'd180     : sin_dat = 16'b0111001000001100 ;  
    10'd181     : sin_dat = 16'b0111001001100101 ;  
    10'd182     : sin_dat = 16'b0111001010111110 ;  
    10'd183     : sin_dat = 16'b0111001100010101 ;  
    10'd184     : sin_dat = 16'b0111001101101011 ;  
    10'd185     : sin_dat = 16'b0111001111000001 ;  
    10'd186     : sin_dat = 16'b0111010000010101 ;  
    10'd187     : sin_dat = 16'b0111010001100111 ;  
    10'd188     : sin_dat = 16'b0111010010111001 ;  
    10'd189     : sin_dat = 16'b0111010100001010 ;  
    10'd190     : sin_dat = 16'b0111010101011001 ;  
    10'd191     : sin_dat = 16'b0111010110101000 ;  
    10'd192     : sin_dat = 16'b0111010111110101 ;  
    10'd193     : sin_dat = 16'b0111011001000001 ;  
    10'd194     : sin_dat = 16'b0111011010001100 ;  
    10'd195     : sin_dat = 16'b0111011011010110 ;  
    10'd196     : sin_dat = 16'b0111011100011110 ;  
    10'd197     : sin_dat = 16'b0111011101100110 ;  
    10'd198     : sin_dat = 16'b0111011110101100 ;  
    10'd199     : sin_dat = 16'b0111011111110010 ;  
    10'd200     : sin_dat = 16'b0111100000110110 ;  
    10'd201     : sin_dat = 16'b0111100001111001 ;  
    10'd202     : sin_dat = 16'b0111100010111010 ;  
    10'd203     : sin_dat = 16'b0111100011111011 ;  
    10'd204     : sin_dat = 16'b0111100100111010 ;  
    10'd205     : sin_dat = 16'b0111100101111000 ;  
    10'd206     : sin_dat = 16'b0111100110110101 ;  
    10'd207     : sin_dat = 16'b0111100111110001 ;  
    10'd208     : sin_dat = 16'b0111101000101100 ;  
    10'd209     : sin_dat = 16'b0111101001100110 ;  
    10'd210     : sin_dat = 16'b0111101010011110 ;  
    10'd211     : sin_dat = 16'b0111101011010101 ;  
    10'd212     : sin_dat = 16'b0111101100001011 ;  
    10'd213     : sin_dat = 16'b0111101101000000 ;  
    10'd214     : sin_dat = 16'b0111101101110011 ;  
    10'd215     : sin_dat = 16'b0111101110100110 ;  
    10'd216     : sin_dat = 16'b0111101111010111 ;  
    10'd217     : sin_dat = 16'b0111110000000111 ;  
    10'd218     : sin_dat = 16'b0111110000110110 ;  
    10'd219     : sin_dat = 16'b0111110001100100 ;  
    10'd220     : sin_dat = 16'b0111110010010000 ;  
    10'd221     : sin_dat = 16'b0111110010111011 ;  
    10'd222     : sin_dat = 16'b0111110011100101 ;  
    10'd223     : sin_dat = 16'b0111110100001110 ;  
    10'd224     : sin_dat = 16'b0111110100110110 ;  
    10'd225     : sin_dat = 16'b0111110101011100 ;  
    10'd226     : sin_dat = 16'b0111110110000001 ;  
    10'd227     : sin_dat = 16'b0111110110100101 ;  
    10'd228     : sin_dat = 16'b0111110111001000 ;  
    10'd229     : sin_dat = 16'b0111110111101010 ;  
    10'd230     : sin_dat = 16'b0111111000001010 ;  
    10'd231     : sin_dat = 16'b0111111000101001 ;  
    10'd232     : sin_dat = 16'b0111111001000111 ;  
    10'd233     : sin_dat = 16'b0111111001100100 ;  
    10'd234     : sin_dat = 16'b0111111001111111 ;  
    10'd235     : sin_dat = 16'b0111111010011001 ;  
    10'd236     : sin_dat = 16'b0111111010110010 ;  
    10'd237     : sin_dat = 16'b0111111011001010 ;  
    10'd238     : sin_dat = 16'b0111111011100001 ;  
    10'd239     : sin_dat = 16'b0111111011110110 ;  
    10'd240     : sin_dat = 16'b0111111100001010 ;  
    10'd241     : sin_dat = 16'b0111111100011101 ;  
    10'd242     : sin_dat = 16'b0111111100101111 ;  
    10'd243     : sin_dat = 16'b0111111100111111 ;  
    10'd244     : sin_dat = 16'b0111111101001111 ;  
    10'd245     : sin_dat = 16'b0111111101011101 ;  
    10'd246     : sin_dat = 16'b0111111101101001 ;  
    10'd247     : sin_dat = 16'b0111111101110101 ;  
    10'd248     : sin_dat = 16'b0111111101111111 ;  
    10'd249     : sin_dat = 16'b0111111110001000 ;  
    10'd250     : sin_dat = 16'b0111111110010000 ;  
    10'd251     : sin_dat = 16'b0111111110010111 ;  
    10'd252     : sin_dat = 16'b0111111110011100 ;  
    10'd253     : sin_dat = 16'b0111111110100000 ;  
    10'd254     : sin_dat = 16'b0111111110100011 ;  
    10'd255     : sin_dat = 16'b0111111110100101 ;  
    10'd256     : sin_dat = 16'b0111111110100101 ;  
    10'd257     : sin_dat = 16'b0111111110100101 ;  
    10'd258     : sin_dat = 16'b0111111110100011 ;  
    10'd259     : sin_dat = 16'b0111111110100000 ;  
    10'd260     : sin_dat = 16'b0111111110011011 ;  
    10'd261     : sin_dat = 16'b0111111110010101 ;  
    10'd262     : sin_dat = 16'b0111111110001110 ;  
    10'd263     : sin_dat = 16'b0111111110000110 ;  
    10'd264     : sin_dat = 16'b0111111101111101 ;  
    10'd265     : sin_dat = 16'b0111111101110010 ;  
    10'd266     : sin_dat = 16'b0111111101100110 ;  
    10'd267     : sin_dat = 16'b0111111101011001 ;  
    10'd268     : sin_dat = 16'b0111111101001011 ;  
    10'd269     : sin_dat = 16'b0111111100111100 ;  
    10'd270     : sin_dat = 16'b0111111100101011 ;  
    10'd271     : sin_dat = 16'b0111111100011001 ;  
    10'd272     : sin_dat = 16'b0111111100000110 ;  
    10'd273     : sin_dat = 16'b0111111011110001 ;  
    10'd274     : sin_dat = 16'b0111111011011100 ;  
    10'd275     : sin_dat = 16'b0111111011000101 ;  
    10'd276     : sin_dat = 16'b0111111010101101 ;  
    10'd277     : sin_dat = 16'b0111111010010011 ;  
    10'd278     : sin_dat = 16'b0111111001111001 ;  
    10'd279     : sin_dat = 16'b0111111001011101 ;  
    10'd280     : sin_dat = 16'b0111111001000000 ;  
    10'd281     : sin_dat = 16'b0111111000100010 ;  
    10'd282     : sin_dat = 16'b0111111000000010 ;  
    10'd283     : sin_dat = 16'b0111110111100010 ;  
    10'd284     : sin_dat = 16'b0111110111000000 ;  
    10'd285     : sin_dat = 16'b0111110110011101 ;  
    10'd286     : sin_dat = 16'b0111110101111000 ;  
    10'd287     : sin_dat = 16'b0111110101010011 ;  
    10'd288     : sin_dat = 16'b0111110100101100 ;  
    10'd289     : sin_dat = 16'b0111110100000100 ;  
    10'd290     : sin_dat = 16'b0111110011011011 ;  
    10'd291     : sin_dat = 16'b0111110010110001 ;  
    10'd292     : sin_dat = 16'b0111110010000101 ;  
    10'd293     : sin_dat = 16'b0111110001011001 ;  
    10'd294     : sin_dat = 16'b0111110000101011 ;  
    10'd295     : sin_dat = 16'b0111101111111100 ;  
    10'd296     : sin_dat = 16'b0111101111001011 ;  
    10'd297     : sin_dat = 16'b0111101110011010 ;  
    10'd298     : sin_dat = 16'b0111101101100111 ;  
    10'd299     : sin_dat = 16'b0111101100110011 ;  
    10'd300     : sin_dat = 16'b0111101011111110 ;  
    10'd301     : sin_dat = 16'b0111101011001000 ;  
    10'd302     : sin_dat = 16'b0111101010010001 ;  
    10'd303     : sin_dat = 16'b0111101001011000 ;  
    10'd304     : sin_dat = 16'b0111101000011110 ;  
    10'd305     : sin_dat = 16'b0111100111100011 ;  
    10'd306     : sin_dat = 16'b0111100110100111 ;  
    10'd307     : sin_dat = 16'b0111100101101010 ;  
    10'd308     : sin_dat = 16'b0111100100101011 ;  
    10'd309     : sin_dat = 16'b0111100011101011 ;  
    10'd310     : sin_dat = 16'b0111100010101011 ;  
    10'd311     : sin_dat = 16'b0111100001101001 ;  
    10'd312     : sin_dat = 16'b0111100000100101 ;  
    10'd313     : sin_dat = 16'b0111011111100001 ;  
    10'd314     : sin_dat = 16'b0111011110011100 ;  
    10'd315     : sin_dat = 16'b0111011101010101 ;  
    10'd316     : sin_dat = 16'b0111011100001101 ;  
    10'd317     : sin_dat = 16'b0111011011000100 ;  
    10'd318     : sin_dat = 16'b0111011001111010 ;  
    10'd319     : sin_dat = 16'b0111011000101111 ;  
    10'd320     : sin_dat = 16'b0111010111100010 ;  
    10'd321     : sin_dat = 16'b0111010110010101 ;  
    10'd322     : sin_dat = 16'b0111010101000110 ;  
    10'd323     : sin_dat = 16'b0111010011110111 ;  
    10'd324     : sin_dat = 16'b0111010010100110 ;  
    10'd325     : sin_dat = 16'b0111010001010100 ;  
    10'd326     : sin_dat = 16'b0111010000000000 ;  
    10'd327     : sin_dat = 16'b0111001110101100 ;  
    10'd328     : sin_dat = 16'b0111001101010111 ;  
    10'd329     : sin_dat = 16'b0111001100000000 ;  
    10'd330     : sin_dat = 16'b0111001010101001 ;  
    10'd331     : sin_dat = 16'b0111001001010000 ;  
    10'd332     : sin_dat = 16'b0111000111110110 ;  
    10'd333     : sin_dat = 16'b0111000110011011 ;  
    10'd334     : sin_dat = 16'b0111000100111111 ;  
    10'd335     : sin_dat = 16'b0111000011100010 ;  
    10'd336     : sin_dat = 16'b0111000010000100 ;  
    10'd337     : sin_dat = 16'b0111000000100101 ;  
    10'd338     : sin_dat = 16'b0110111111000100 ;  
    10'd339     : sin_dat = 16'b0110111101100011 ;  
    10'd340     : sin_dat = 16'b0110111100000000 ;  
    10'd341     : sin_dat = 16'b0110111010011101 ;  
    10'd342     : sin_dat = 16'b0110111000111000 ;  
    10'd343     : sin_dat = 16'b0110110111010010 ;  
    10'd344     : sin_dat = 16'b0110110101101100 ;  
    10'd345     : sin_dat = 16'b0110110100000100 ;  
    10'd346     : sin_dat = 16'b0110110010011011 ;  
    10'd347     : sin_dat = 16'b0110110000110001 ;  
    10'd348     : sin_dat = 16'b0110101111000110 ;  
    10'd349     : sin_dat = 16'b0110101101011010 ;  
    10'd350     : sin_dat = 16'b0110101011101101 ;  
    10'd351     : sin_dat = 16'b0110101001111111 ;  
    10'd352     : sin_dat = 16'b0110101000010000 ;  
    10'd353     : sin_dat = 16'b0110100110100000 ;  
    10'd354     : sin_dat = 16'b0110100100101111 ;  
    10'd355     : sin_dat = 16'b0110100010111100 ;  
    10'd356     : sin_dat = 16'b0110100001001001 ;  
    10'd357     : sin_dat = 16'b0110011111010101 ;  
    10'd358     : sin_dat = 16'b0110011101100000 ;  
    10'd359     : sin_dat = 16'b0110011011101010 ;  
    10'd360     : sin_dat = 16'b0110011001110010 ;  
    10'd361     : sin_dat = 16'b0110010111111010 ;  
    10'd362     : sin_dat = 16'b0110010110000001 ;  
    10'd363     : sin_dat = 16'b0110010100000111 ;  
    10'd364     : sin_dat = 16'b0110010010001100 ;  
    10'd365     : sin_dat = 16'b0110010000010000 ;  
    10'd366     : sin_dat = 16'b0110001110010011 ;  
    10'd367     : sin_dat = 16'b0110001100010101 ;  
    10'd368     : sin_dat = 16'b0110001010010110 ;  
    10'd369     : sin_dat = 16'b0110001000010110 ;  
    10'd370     : sin_dat = 16'b0110000110010101 ;  
    10'd371     : sin_dat = 16'b0110000100010011 ;  
    10'd372     : sin_dat = 16'b0110000010010001 ;  
    10'd373     : sin_dat = 16'b0110000000001101 ;  
    10'd374     : sin_dat = 16'b0101111110001000 ;  
    10'd375     : sin_dat = 16'b0101111100000011 ;  
    10'd376     : sin_dat = 16'b0101111001111100 ;  
    10'd377     : sin_dat = 16'b0101110111110101 ;  
    10'd378     : sin_dat = 16'b0101110101101101 ;  
    10'd379     : sin_dat = 16'b0101110011100100 ;  
    10'd380     : sin_dat = 16'b0101110001011010 ;  
    10'd381     : sin_dat = 16'b0101101111001111 ;  
    10'd382     : sin_dat = 16'b0101101101000011 ;  
    10'd383     : sin_dat = 16'b0101101010110110 ;  
    10'd384     : sin_dat = 16'b0101101000101001 ;  
    10'd385     : sin_dat = 16'b0101100110011010 ;  
    10'd386     : sin_dat = 16'b0101100100001011 ;  
    10'd387     : sin_dat = 16'b0101100001111011 ;  
    10'd388     : sin_dat = 16'b0101011111101010 ;  
    10'd389     : sin_dat = 16'b0101011101011000 ;  
    10'd390     : sin_dat = 16'b0101011011000101 ;  
    10'd391     : sin_dat = 16'b0101011000110010 ;  
    10'd392     : sin_dat = 16'b0101010110011101 ;  
    10'd393     : sin_dat = 16'b0101010100001000 ;  
    10'd394     : sin_dat = 16'b0101010001110010 ;  
    10'd395     : sin_dat = 16'b0101001111011011 ;  
    10'd396     : sin_dat = 16'b0101001101000100 ;  
    10'd397     : sin_dat = 16'b0101001010101011 ;  
    10'd398     : sin_dat = 16'b0101001000010010 ;  
    10'd399     : sin_dat = 16'b0101000101111000 ;  
    10'd400     : sin_dat = 16'b0101000011011101 ;  
    10'd401     : sin_dat = 16'b0101000001000001 ;  
    10'd402     : sin_dat = 16'b0100111110100101 ;  
    10'd403     : sin_dat = 16'b0100111100001000 ;  
    10'd404     : sin_dat = 16'b0100111001101010 ;  
    10'd405     : sin_dat = 16'b0100110111001011 ;  
    10'd406     : sin_dat = 16'b0100110100101100 ;  
    10'd407     : sin_dat = 16'b0100110010001100 ;  
    10'd408     : sin_dat = 16'b0100101111101011 ;  
    10'd409     : sin_dat = 16'b0100101101001001 ;  
    10'd410     : sin_dat = 16'b0100101010100111 ;  
    10'd411     : sin_dat = 16'b0100101000000100 ;  
    10'd412     : sin_dat = 16'b0100100101100000 ;  
    10'd413     : sin_dat = 16'b0100100010111011 ;  
    10'd414     : sin_dat = 16'b0100100000010110 ;  
    10'd415     : sin_dat = 16'b0100011101110000 ;  
    10'd416     : sin_dat = 16'b0100011011001010 ;  
    10'd417     : sin_dat = 16'b0100011000100011 ;  
    10'd418     : sin_dat = 16'b0100010101111011 ;  
    10'd419     : sin_dat = 16'b0100010011010010 ;  
    10'd420     : sin_dat = 16'b0100010000101001 ;  
    10'd421     : sin_dat = 16'b0100001101111111 ;  
    10'd422     : sin_dat = 16'b0100001011010100 ;  
    10'd423     : sin_dat = 16'b0100001000101001 ;  
    10'd424     : sin_dat = 16'b0100000101111101 ;  
    10'd425     : sin_dat = 16'b0100000011010001 ;  
    10'd426     : sin_dat = 16'b0100000000100011 ;  
    10'd427     : sin_dat = 16'b0011111101110110 ;  
    10'd428     : sin_dat = 16'b0011111011000111 ;  
    10'd429     : sin_dat = 16'b0011111000011000 ;  
    10'd430     : sin_dat = 16'b0011110101101001 ;  
    10'd431     : sin_dat = 16'b0011110010111001 ;  
    10'd432     : sin_dat = 16'b0011110000001000 ;  
    10'd433     : sin_dat = 16'b0011101101010111 ;  
    10'd434     : sin_dat = 16'b0011101010100101 ;  
    10'd435     : sin_dat = 16'b0011100111110010 ;  
    10'd436     : sin_dat = 16'b0011100100111111 ;  
    10'd437     : sin_dat = 16'b0011100010001100 ;  
    10'd438     : sin_dat = 16'b0011011111010111 ;  
    10'd439     : sin_dat = 16'b0011011100100011 ;  
    10'd440     : sin_dat = 16'b0011011001101110 ;  
    10'd441     : sin_dat = 16'b0011010110111000 ;  
    10'd442     : sin_dat = 16'b0011010100000010 ;  
    10'd443     : sin_dat = 16'b0011010001001011 ;  
    10'd444     : sin_dat = 16'b0011001110010100 ;  
    10'd445     : sin_dat = 16'b0011001011011100 ;  
    10'd446     : sin_dat = 16'b0011001000100100 ;  
    10'd447     : sin_dat = 16'b0011000101101011 ;  
    10'd448     : sin_dat = 16'b0011000010110010 ;  
    10'd449     : sin_dat = 16'b0010111111111000 ;  
    10'd450     : sin_dat = 16'b0010111100111110 ;  
    10'd451     : sin_dat = 16'b0010111010000011 ;  
    10'd452     : sin_dat = 16'b0010110111001000 ;  
    10'd453     : sin_dat = 16'b0010110100001101 ;  
    10'd454     : sin_dat = 16'b0010110001010001 ;  
    10'd455     : sin_dat = 16'b0010101110010101 ;  
    10'd456     : sin_dat = 16'b0010101011011000 ;  
    10'd457     : sin_dat = 16'b0010101000011011 ;  
    10'd458     : sin_dat = 16'b0010100101011101 ;  
    10'd459     : sin_dat = 16'b0010100010011111 ;  
    10'd460     : sin_dat = 16'b0010011111100001 ;  
    10'd461     : sin_dat = 16'b0010011100100010 ;  
    10'd462     : sin_dat = 16'b0010011001100011 ;  
    10'd463     : sin_dat = 16'b0010010110100011 ;  
    10'd464     : sin_dat = 16'b0010010011100100 ;  
    10'd465     : sin_dat = 16'b0010010000100011 ;  
    10'd466     : sin_dat = 16'b0010001101100011 ;  
    10'd467     : sin_dat = 16'b0010001010100010 ;  
    10'd468     : sin_dat = 16'b0010000111100001 ;  
    10'd469     : sin_dat = 16'b0010000100011111 ;  
    10'd470     : sin_dat = 16'b0010000001011101 ;  
    10'd471     : sin_dat = 16'b0001111110011011 ;  
    10'd472     : sin_dat = 16'b0001111011011000 ;  
    10'd473     : sin_dat = 16'b0001111000010110 ;  
    10'd474     : sin_dat = 16'b0001110101010011 ;  
    10'd475     : sin_dat = 16'b0001110010001111 ;  
    10'd476     : sin_dat = 16'b0001101111001100 ;  
    10'd477     : sin_dat = 16'b0001101100001000 ;  
    10'd478     : sin_dat = 16'b0001101001000011 ;  
    10'd479     : sin_dat = 16'b0001100101111111 ;  
    10'd480     : sin_dat = 16'b0001100010111010 ;  
    10'd481     : sin_dat = 16'b0001011111110101 ;  
    10'd482     : sin_dat = 16'b0001011100110000 ;  
    10'd483     : sin_dat = 16'b0001011001101011 ;  
    10'd484     : sin_dat = 16'b0001010110100101 ;  
    10'd485     : sin_dat = 16'b0001010011011111 ;  
    10'd486     : sin_dat = 16'b0001010000011001 ;  
    10'd487     : sin_dat = 16'b0001001101010011 ;  
    10'd488     : sin_dat = 16'b0001001010001101 ;  
    10'd489     : sin_dat = 16'b0001000111000110 ;  
    10'd490     : sin_dat = 16'b0001000100000000 ;  
    10'd491     : sin_dat = 16'b0001000000111001 ;  
    10'd492     : sin_dat = 16'b0000111101110010 ;  
    10'd493     : sin_dat = 16'b0000111010101010 ;  
    10'd494     : sin_dat = 16'b0000110111100011 ;  
    10'd495     : sin_dat = 16'b0000110100011100 ;  
    10'd496     : sin_dat = 16'b0000110001010100 ;  
    10'd497     : sin_dat = 16'b0000101110001100 ;  
    10'd498     : sin_dat = 16'b0000101011000100 ;  
    10'd499     : sin_dat = 16'b0000100111111100 ;  
    10'd500     : sin_dat = 16'b0000100100110100 ;  
    10'd501     : sin_dat = 16'b0000100001101100 ;  
    10'd502     : sin_dat = 16'b0000011110100100 ;  
    10'd503     : sin_dat = 16'b0000011011011100 ;  
    10'd504     : sin_dat = 16'b0000011000010011 ;  
    10'd505     : sin_dat = 16'b0000010101001011 ;  
    10'd506     : sin_dat = 16'b0000010010000011 ;  
    10'd507     : sin_dat = 16'b0000001110111010 ;  
    10'd508     : sin_dat = 16'b0000001011110010 ;  
    10'd509     : sin_dat = 16'b0000001000101001 ;  
    10'd510     : sin_dat = 16'b0000000101100000 ;  
    10'd511     : sin_dat = 16'b0000000010011000 ;  
    10'd512     : sin_dat = 16'b1111111111001111 ;  
    10'd513     : sin_dat = 16'b1111111100000111 ;  
    10'd514     : sin_dat = 16'b1111111000111110 ;  
    10'd515     : sin_dat = 16'b1111110101110101 ;  
    10'd516     : sin_dat = 16'b1111110010101101 ;  
    10'd517     : sin_dat = 16'b1111101111100100 ;  
    10'd518     : sin_dat = 16'b1111101100011100 ;  
    10'd519     : sin_dat = 16'b1111101001010011 ;  
    10'd520     : sin_dat = 16'b1111100110001011 ;  
    10'd521     : sin_dat = 16'b1111100011000011 ;  
    10'd522     : sin_dat = 16'b1111011111111011 ;  
    10'd523     : sin_dat = 16'b1111011100110010 ;  
    10'd524     : sin_dat = 16'b1111011001101010 ;  
    10'd525     : sin_dat = 16'b1111010110100010 ;  
    10'd526     : sin_dat = 16'b1111010011011010 ;  
    10'd527     : sin_dat = 16'b1111010000010011 ;  
    10'd528     : sin_dat = 16'b1111001101001011 ;  
    10'd529     : sin_dat = 16'b1111001010000011 ;  
    10'd530     : sin_dat = 16'b1111000110111100 ;  
    10'd531     : sin_dat = 16'b1111000011110101 ;  
    10'd532     : sin_dat = 16'b1111000000101110 ;  
    10'd533     : sin_dat = 16'b1110111101100111 ;  
    10'd534     : sin_dat = 16'b1110111010100000 ;  
    10'd535     : sin_dat = 16'b1110110111011001 ;  
    10'd536     : sin_dat = 16'b1110110100010011 ;  
    10'd537     : sin_dat = 16'b1110110001001100 ;  
    10'd538     : sin_dat = 16'b1110101110000110 ;  
    10'd539     : sin_dat = 16'b1110101011000000 ;  
    10'd540     : sin_dat = 16'b1110100111111011 ;  
    10'd541     : sin_dat = 16'b1110100100110101 ;  
    10'd542     : sin_dat = 16'b1110100001110000 ;  
    10'd543     : sin_dat = 16'b1110011110101011 ;  
    10'd544     : sin_dat = 16'b1110011011100110 ;  
    10'd545     : sin_dat = 16'b1110011000100001 ;  
    10'd546     : sin_dat = 16'b1110010101011101 ;  
    10'd547     : sin_dat = 16'b1110010010011001 ;  
    10'd548     : sin_dat = 16'b1110001111010101 ;  
    10'd549     : sin_dat = 16'b1110001100010010 ;  
    10'd550     : sin_dat = 16'b1110001001001111 ;  
    10'd551     : sin_dat = 16'b1110000110001100 ;  
    10'd552     : sin_dat = 16'b1110000011001001 ;  
    10'd553     : sin_dat = 16'b1110000000000111 ;  
    10'd554     : sin_dat = 16'b1101111101000101 ;  
    10'd555     : sin_dat = 16'b1101111010000011 ;  
    10'd556     : sin_dat = 16'b1101110111000001 ;  
    10'd557     : sin_dat = 16'b1101110100000000 ;  
    10'd558     : sin_dat = 16'b1101110001000000 ;  
    10'd559     : sin_dat = 16'b1101101101111111 ;  
    10'd560     : sin_dat = 16'b1101101010111111 ;  
    10'd561     : sin_dat = 16'b1101100111111111 ;  
    10'd562     : sin_dat = 16'b1101100101000000 ;  
    10'd563     : sin_dat = 16'b1101100010000001 ;  
    10'd564     : sin_dat = 16'b1101011111000011 ;  
    10'd565     : sin_dat = 16'b1101011100000100 ;  
    10'd566     : sin_dat = 16'b1101011001000111 ;  
    10'd567     : sin_dat = 16'b1101010110001001 ;  
    10'd568     : sin_dat = 16'b1101010011001100 ;  
    10'd569     : sin_dat = 16'b1101010000010000 ;  
    10'd570     : sin_dat = 16'b1101001101010100 ;  
    10'd571     : sin_dat = 16'b1101001010011000 ;  
    10'd572     : sin_dat = 16'b1101000111011101 ;  
    10'd573     : sin_dat = 16'b1101000100100010 ;  
    10'd574     : sin_dat = 16'b1101000001100111 ;  
    10'd575     : sin_dat = 16'b1100111110101101 ;  
    10'd576     : sin_dat = 16'b1100111011110100 ;  
    10'd577     : sin_dat = 16'b1100111000111011 ;  
    10'd578     : sin_dat = 16'b1100110110000011 ;  
    10'd579     : sin_dat = 16'b1100110011001011 ;  
    10'd580     : sin_dat = 16'b1100110000010011 ;  
    10'd581     : sin_dat = 16'b1100101101011100 ;  
    10'd582     : sin_dat = 16'b1100101010100110 ;  
    10'd583     : sin_dat = 16'b1100100111110000 ;  
    10'd584     : sin_dat = 16'b1100100100111010 ;  
    10'd585     : sin_dat = 16'b1100100010000101 ;  
    10'd586     : sin_dat = 16'b1100011111010001 ;  
    10'd587     : sin_dat = 16'b1100011100011101 ;  
    10'd588     : sin_dat = 16'b1100011001101010 ;  
    10'd589     : sin_dat = 16'b1100010110110111 ;  
    10'd590     : sin_dat = 16'b1100010100000101 ;  
    10'd591     : sin_dat = 16'b1100010001010011 ;  
    10'd592     : sin_dat = 16'b1100001110100010 ;  
    10'd593     : sin_dat = 16'b1100001011110010 ;  
    10'd594     : sin_dat = 16'b1100001001000010 ;  
    10'd595     : sin_dat = 16'b1100000110010010 ;  
    10'd596     : sin_dat = 16'b1100000011100100 ;  
    10'd597     : sin_dat = 16'b1100000000110110 ;  
    10'd598     : sin_dat = 16'b1011111110001000 ;  
    10'd599     : sin_dat = 16'b1011111011011011 ;  
    10'd600     : sin_dat = 16'b1011111000101111 ;  
    10'd601     : sin_dat = 16'b1011110110000100 ;  
    10'd602     : sin_dat = 16'b1011110011011001 ;  
    10'd603     : sin_dat = 16'b1011110000101110 ;  
    10'd604     : sin_dat = 16'b1011101110000101 ;  
    10'd605     : sin_dat = 16'b1011101011011100 ;  
    10'd606     : sin_dat = 16'b1011101000110100 ;  
    10'd607     : sin_dat = 16'b1011100110001100 ;  
    10'd608     : sin_dat = 16'b1011100011100101 ;  
    10'd609     : sin_dat = 16'b1011100000111111 ;  
    10'd610     : sin_dat = 16'b1011011110011001 ;  
    10'd611     : sin_dat = 16'b1011011011110100 ;  
    10'd612     : sin_dat = 16'b1011011001010000 ;  
    10'd613     : sin_dat = 16'b1011010110101101 ;  
    10'd614     : sin_dat = 16'b1011010100001010 ;  
    10'd615     : sin_dat = 16'b1011010001101000 ;  
    10'd616     : sin_dat = 16'b1011001111000111 ;  
    10'd617     : sin_dat = 16'b1011001100100110 ;  
    10'd618     : sin_dat = 16'b1011001010000110 ;  
    10'd619     : sin_dat = 16'b1011000111100111 ;  
    10'd620     : sin_dat = 16'b1011000101001001 ;  
    10'd621     : sin_dat = 16'b1011000010101011 ;  
    10'd622     : sin_dat = 16'b1011000000001111 ;  
    10'd623     : sin_dat = 16'b1010111101110011 ;  
    10'd624     : sin_dat = 16'b1010111011010111 ;  
    10'd625     : sin_dat = 16'b1010111000111101 ;  
    10'd626     : sin_dat = 16'b1010110110100011 ;  
    10'd627     : sin_dat = 16'b1010110100001010 ;  
    10'd628     : sin_dat = 16'b1010110001110010 ;  
    10'd629     : sin_dat = 16'b1010101111011011 ;  
    10'd630     : sin_dat = 16'b1010101101000101 ;  
    10'd631     : sin_dat = 16'b1010101010101111 ;  
    10'd632     : sin_dat = 16'b1010101000011010 ;  
    10'd633     : sin_dat = 16'b1010100110000110 ;  
    10'd634     : sin_dat = 16'b1010100011110011 ;  
    10'd635     : sin_dat = 16'b1010100001100001 ;  
    10'd636     : sin_dat = 16'b1010011111001111 ;  
    10'd637     : sin_dat = 16'b1010011100111111 ;  
    10'd638     : sin_dat = 16'b1010011010101111 ;  
    10'd639     : sin_dat = 16'b1010011000100000 ;  
    10'd640     : sin_dat = 16'b1010010110010010 ;  
    10'd641     : sin_dat = 16'b1010010100000101 ;  
    10'd642     : sin_dat = 16'b1010010001111001 ;  
    10'd643     : sin_dat = 16'b1010001111101101 ;  
    10'd644     : sin_dat = 16'b1010001101100011 ;  
    10'd645     : sin_dat = 16'b1010001011011001 ;  
    10'd646     : sin_dat = 16'b1010001001010000 ;  
    10'd647     : sin_dat = 16'b1010000111001001 ;  
    10'd648     : sin_dat = 16'b1010000101000010 ;  
    10'd649     : sin_dat = 16'b1010000010111100 ;  
    10'd650     : sin_dat = 16'b1010000000110111 ;  
    10'd651     : sin_dat = 16'b1001111110110011 ;  
    10'd652     : sin_dat = 16'b1001111100101111 ;  
    10'd653     : sin_dat = 16'b1001111010101101 ;  
    10'd654     : sin_dat = 16'b1001111000101100 ;  
    10'd655     : sin_dat = 16'b1001110110101011 ;  
    10'd656     : sin_dat = 16'b1001110100101100 ;  
    10'd657     : sin_dat = 16'b1001110010101101 ;  
    10'd658     : sin_dat = 16'b1001110000110000 ;  
    10'd659     : sin_dat = 16'b1001101110110011 ;  
    10'd660     : sin_dat = 16'b1001101100111000 ;  
    10'd661     : sin_dat = 16'b1001101010111101 ;  
    10'd662     : sin_dat = 16'b1001101001000011 ;  
    10'd663     : sin_dat = 16'b1001100111001011 ;  
    10'd664     : sin_dat = 16'b1001100101010011 ;  
    10'd665     : sin_dat = 16'b1001100011011100 ;  
    10'd666     : sin_dat = 16'b1001100001100111 ;  
    10'd667     : sin_dat = 16'b1001011111110010 ;  
    10'd668     : sin_dat = 16'b1001011101111110 ;  
    10'd669     : sin_dat = 16'b1001011100001100 ;  
    10'd670     : sin_dat = 16'b1001011010011010 ;  
    10'd671     : sin_dat = 16'b1001011000101001 ;  
    10'd672     : sin_dat = 16'b1001010110111010 ;  
    10'd673     : sin_dat = 16'b1001010101001011 ;  
    10'd674     : sin_dat = 16'b1001010011011101 ;  
    10'd675     : sin_dat = 16'b1001010001110001 ;  
    10'd676     : sin_dat = 16'b1001010000000101 ;  
    10'd677     : sin_dat = 16'b1001001110011011 ;  
    10'd678     : sin_dat = 16'b1001001100110001 ;  
    10'd679     : sin_dat = 16'b1001001011001001 ;  
    10'd680     : sin_dat = 16'b1001001001100010 ;  
    10'd681     : sin_dat = 16'b1001000111111011 ;  
    10'd682     : sin_dat = 16'b1001000110010110 ;  
    10'd683     : sin_dat = 16'b1001000100110010 ;  
    10'd684     : sin_dat = 16'b1001000011001111 ;  
    10'd685     : sin_dat = 16'b1001000001101101 ;  
    10'd686     : sin_dat = 16'b1001000000001100 ;  
    10'd687     : sin_dat = 16'b1000111110101100 ;  
    10'd688     : sin_dat = 16'b1000111101001110 ;  
    10'd689     : sin_dat = 16'b1000111011110000 ;  
    10'd690     : sin_dat = 16'b1000111010010011 ;  
    10'd691     : sin_dat = 16'b1000111000111000 ;  
    10'd692     : sin_dat = 16'b1000110111011101 ;  
    10'd693     : sin_dat = 16'b1000110110000100 ;  
    10'd694     : sin_dat = 16'b1000110100101100 ;  
    10'd695     : sin_dat = 16'b1000110011010101 ;  
    10'd696     : sin_dat = 16'b1000110001111111 ;  
    10'd697     : sin_dat = 16'b1000110000101010 ;  
    10'd698     : sin_dat = 16'b1000101111010110 ;  
    10'd699     : sin_dat = 16'b1000101110000100 ;  
    10'd700     : sin_dat = 16'b1000101100110010 ;  
    10'd701     : sin_dat = 16'b1000101011100010 ;  
    10'd702     : sin_dat = 16'b1000101010010011 ;  
    10'd703     : sin_dat = 16'b1000101001000101 ;  
    10'd704     : sin_dat = 16'b1000100111111000 ;  
    10'd705     : sin_dat = 16'b1000100110101100 ;  
    10'd706     : sin_dat = 16'b1000100101100001 ;  
    10'd707     : sin_dat = 16'b1000100100011000 ;  
    10'd708     : sin_dat = 16'b1000100011001111 ;  
    10'd709     : sin_dat = 16'b1000100010001000 ;  
    10'd710     : sin_dat = 16'b1000100001000010 ;  
    10'd711     : sin_dat = 16'b1000011111111101 ;  
    10'd712     : sin_dat = 16'b1000011110111001 ;  
    10'd713     : sin_dat = 16'b1000011101110111 ;  
    10'd714     : sin_dat = 16'b1000011100110101 ;  
    10'd715     : sin_dat = 16'b1000011011110101 ;  
    10'd716     : sin_dat = 16'b1000011010110110 ;  
    10'd717     : sin_dat = 16'b1000011001111000 ;  
    10'd718     : sin_dat = 16'b1000011000111011 ;  
    10'd719     : sin_dat = 16'b1000010111111111 ;  
    10'd720     : sin_dat = 16'b1000010111000101 ;  
    10'd721     : sin_dat = 16'b1000010110001100 ;  
    10'd722     : sin_dat = 16'b1000010101010100 ;  
    10'd723     : sin_dat = 16'b1000010100011101 ;  
    10'd724     : sin_dat = 16'b1000010011100111 ;  
    10'd725     : sin_dat = 16'b1000010010110011 ;  
    10'd726     : sin_dat = 16'b1000010001111111 ;  
    10'd727     : sin_dat = 16'b1000010001001101 ;  
    10'd728     : sin_dat = 16'b1000010000011100 ;  
    10'd729     : sin_dat = 16'b1000001111101100 ;  
    10'd730     : sin_dat = 16'b1000001110111110 ;  
    10'd731     : sin_dat = 16'b1000001110010001 ;  
    10'd732     : sin_dat = 16'b1000001101100100 ;  
    10'd733     : sin_dat = 16'b1000001100111010 ;  
    10'd734     : sin_dat = 16'b1000001100010000 ;  
    10'd735     : sin_dat = 16'b1000001011100111 ;  
    10'd736     : sin_dat = 16'b1000001011000000 ;  
    10'd737     : sin_dat = 16'b1000001010011010 ;  
    10'd738     : sin_dat = 16'b1000001001110101 ;  
    10'd739     : sin_dat = 16'b1000001001010001 ;  
    10'd740     : sin_dat = 16'b1000001000101111 ;  
    10'd741     : sin_dat = 16'b1000001000001101 ;  
    10'd742     : sin_dat = 16'b1000000111101101 ;  
    10'd743     : sin_dat = 16'b1000000111001111 ;  
    10'd744     : sin_dat = 16'b1000000110110001 ;  
    10'd745     : sin_dat = 16'b1000000110010101 ;  
    10'd746     : sin_dat = 16'b1000000101111001 ;  
    10'd747     : sin_dat = 16'b1000000101011111 ;  
    10'd748     : sin_dat = 16'b1000000101000111 ;  
    10'd749     : sin_dat = 16'b1000000100101111 ;  
    10'd750     : sin_dat = 16'b1000000100011001 ;  
    10'd751     : sin_dat = 16'b1000000100000100 ;  
    10'd752     : sin_dat = 16'b1000000011110000 ;  
    10'd753     : sin_dat = 16'b1000000011011101 ;  
    10'd754     : sin_dat = 16'b1000000011001100 ;  
    10'd755     : sin_dat = 16'b1000000010111100 ;  
    10'd756     : sin_dat = 16'b1000000010101101 ;  
    10'd757     : sin_dat = 16'b1000000010011111 ;  
    10'd758     : sin_dat = 16'b1000000010010011 ;  
    10'd759     : sin_dat = 16'b1000000010000111 ;  
    10'd760     : sin_dat = 16'b1000000001111101 ;  
    10'd761     : sin_dat = 16'b1000000001110101 ;  
    10'd762     : sin_dat = 16'b1000000001101101 ;  
    10'd763     : sin_dat = 16'b1000000001100111 ;  
    10'd764     : sin_dat = 16'b1000000001100010 ;  
    10'd765     : sin_dat = 16'b1000000001011110 ;  
    10'd766     : sin_dat = 16'b1000000001011011 ;  
    10'd767     : sin_dat = 16'b1000000001011010 ;  
    10'd768     : sin_dat = 16'b1000000001011010 ;  
    10'd769     : sin_dat = 16'b1000000001011011 ;  
    10'd770     : sin_dat = 16'b1000000001011101 ;  
    10'd771     : sin_dat = 16'b1000000001100000 ;  
    10'd772     : sin_dat = 16'b1000000001100101 ;  
    10'd773     : sin_dat = 16'b1000000001101011 ;  
    10'd774     : sin_dat = 16'b1000000001110010 ;  
    10'd775     : sin_dat = 16'b1000000001111011 ;  
    10'd776     : sin_dat = 16'b1000000010000101 ;  
    10'd777     : sin_dat = 16'b1000000010001111 ;  
    10'd778     : sin_dat = 16'b1000000010011100 ;  
    10'd779     : sin_dat = 16'b1000000010101001 ;  
    10'd780     : sin_dat = 16'b1000000010111000 ;  
    10'd781     : sin_dat = 16'b1000000011000111 ;  
    10'd782     : sin_dat = 16'b1000000011011000 ;  
    10'd783     : sin_dat = 16'b1000000011101011 ;  
    10'd784     : sin_dat = 16'b1000000011111110 ;  
    10'd785     : sin_dat = 16'b1000000100010011 ;  
    10'd786     : sin_dat = 16'b1000000100101001 ;  
    10'd787     : sin_dat = 16'b1000000101000000 ;  
    10'd788     : sin_dat = 16'b1000000101011000 ;  
    10'd789     : sin_dat = 16'b1000000101110010 ;  
    10'd790     : sin_dat = 16'b1000000110001101 ;  
    10'd791     : sin_dat = 16'b1000000110101001 ;  
    10'd792     : sin_dat = 16'b1000000111000110 ;  
    10'd793     : sin_dat = 16'b1000000111100101 ;  
    10'd794     : sin_dat = 16'b1000001000000100 ;  
    10'd795     : sin_dat = 16'b1000001000100101 ;  
    10'd796     : sin_dat = 16'b1000001001001000 ;  
    10'd797     : sin_dat = 16'b1000001001101011 ;  
    10'd798     : sin_dat = 16'b1000001010001111 ;  
    10'd799     : sin_dat = 16'b1000001010110101 ;  
    10'd800     : sin_dat = 16'b1000001011011100 ;  
    10'd801     : sin_dat = 16'b1000001100000100 ;  
    10'd802     : sin_dat = 16'b1000001100101110 ;  
    10'd803     : sin_dat = 16'b1000001101011000 ;  
    10'd804     : sin_dat = 16'b1000001110000100 ;  
    10'd805     : sin_dat = 16'b1000001110110001 ;  
    10'd806     : sin_dat = 16'b1000001111011111 ;  
    10'd807     : sin_dat = 16'b1000010000001111 ;  
    10'd808     : sin_dat = 16'b1000010000111111 ;  
    10'd809     : sin_dat = 16'b1000010001110001 ;  
    10'd810     : sin_dat = 16'b1000010010100100 ;  
    10'd811     : sin_dat = 16'b1000010011011000 ;  
    10'd812     : sin_dat = 16'b1000010100001110 ;  
    10'd813     : sin_dat = 16'b1000010101000100 ;  
    10'd814     : sin_dat = 16'b1000010101111100 ;  
    10'd815     : sin_dat = 16'b1000010110110101 ;  
    10'd816     : sin_dat = 16'b1000010111101111 ;  
    10'd817     : sin_dat = 16'b1000011000101010 ;  
    10'd818     : sin_dat = 16'b1000011001100111 ;  
    10'd819     : sin_dat = 16'b1000011010100100 ;  
    10'd820     : sin_dat = 16'b1000011011100011 ;  
    10'd821     : sin_dat = 16'b1000011100100011 ;  
    10'd822     : sin_dat = 16'b1000011101100100 ;  
    10'd823     : sin_dat = 16'b1000011110100111 ;  
    10'd824     : sin_dat = 16'b1000011111101010 ;  
    10'd825     : sin_dat = 16'b1000100000101111 ;  
    10'd826     : sin_dat = 16'b1000100001110100 ;  
    10'd827     : sin_dat = 16'b1000100010111011 ;  
    10'd828     : sin_dat = 16'b1000100100000011 ;  
    10'd829     : sin_dat = 16'b1000100101001101 ;  
    10'd830     : sin_dat = 16'b1000100110010111 ;  
    10'd831     : sin_dat = 16'b1000100111100010 ;  
    10'd832     : sin_dat = 16'b1000101000101111 ;  
    10'd833     : sin_dat = 16'b1000101001111101 ;  
    10'd834     : sin_dat = 16'b1000101011001100 ;  
    10'd835     : sin_dat = 16'b1000101100011100 ;  
    10'd836     : sin_dat = 16'b1000101101101101 ;  
    10'd837     : sin_dat = 16'b1000101110111111 ;  
    10'd838     : sin_dat = 16'b1000110000010011 ;  
    10'd839     : sin_dat = 16'b1000110001100111 ;  
    10'd840     : sin_dat = 16'b1000110010111101 ;  
    10'd841     : sin_dat = 16'b1000110100010100 ;  
    10'd842     : sin_dat = 16'b1000110101101100 ;  
    10'd843     : sin_dat = 16'b1000110111000100 ;  
    10'd844     : sin_dat = 16'b1000111000011111 ;  
    10'd845     : sin_dat = 16'b1000111001111010 ;  
    10'd846     : sin_dat = 16'b1000111011010110 ;  
    10'd847     : sin_dat = 16'b1000111100110011 ;  
    10'd848     : sin_dat = 16'b1000111110010010 ;  
    10'd849     : sin_dat = 16'b1000111111110001 ;  
    10'd850     : sin_dat = 16'b1001000001010010 ;  
    10'd851     : sin_dat = 16'b1001000010110100 ;  
    10'd852     : sin_dat = 16'b1001000100010110 ;  
    10'd853     : sin_dat = 16'b1001000101111010 ;  
    10'd854     : sin_dat = 16'b1001000111011111 ;  
    10'd855     : sin_dat = 16'b1001001001000101 ;  
    10'd856     : sin_dat = 16'b1001001010101100 ;  
    10'd857     : sin_dat = 16'b1001001100010100 ;  
    10'd858     : sin_dat = 16'b1001001101111101 ;  
    10'd859     : sin_dat = 16'b1001001111101000 ;  
    10'd860     : sin_dat = 16'b1001010001010011 ;  
    10'd861     : sin_dat = 16'b1001010010111111 ;  
    10'd862     : sin_dat = 16'b1001010100101100 ;  
    10'd863     : sin_dat = 16'b1001010110011011 ;  
    10'd864     : sin_dat = 16'b1001011000001010 ;  
    10'd865     : sin_dat = 16'b1001011001111010 ;  
    10'd866     : sin_dat = 16'b1001011011101100 ;  
    10'd867     : sin_dat = 16'b1001011101011110 ;  
    10'd868     : sin_dat = 16'b1001011111010010 ;  
    10'd869     : sin_dat = 16'b1001100001000110 ;  
    10'd870     : sin_dat = 16'b1001100010111011 ;  
    10'd871     : sin_dat = 16'b1001100100110010 ;  
    10'd872     : sin_dat = 16'b1001100110101001 ;  
    10'd873     : sin_dat = 16'b1001101000100010 ;  
    10'd874     : sin_dat = 16'b1001101010011011 ;  
    10'd875     : sin_dat = 16'b1001101100010101 ;  
    10'd876     : sin_dat = 16'b1001101110010001 ;  
    10'd877     : sin_dat = 16'b1001110000001101 ;  
    10'd878     : sin_dat = 16'b1001110010001010 ;  
    10'd879     : sin_dat = 16'b1001110100001001 ;  
    10'd880     : sin_dat = 16'b1001110110001000 ;  
    10'd881     : sin_dat = 16'b1001111000001000 ;  
    10'd882     : sin_dat = 16'b1001111010001001 ;  
    10'd883     : sin_dat = 16'b1001111100001011 ;  
    10'd884     : sin_dat = 16'b1001111110001110 ;  
    10'd885     : sin_dat = 16'b1010000000010010 ;  
    10'd886     : sin_dat = 16'b1010000010010111 ;  
    10'd887     : sin_dat = 16'b1010000100011100 ;  
    10'd888     : sin_dat = 16'b1010000110100011 ;  
    10'd889     : sin_dat = 16'b1010001000101011 ;  
    10'd890     : sin_dat = 16'b1010001010110011 ;  
    10'd891     : sin_dat = 16'b1010001100111100 ;  
    10'd892     : sin_dat = 16'b1010001111000111 ;  
    10'd893     : sin_dat = 16'b1010010001010010 ;  
    10'd894     : sin_dat = 16'b1010010011011110 ;  
    10'd895     : sin_dat = 16'b1010010101101011 ;  
    10'd896     : sin_dat = 16'b1010010111111000 ;  
    10'd897     : sin_dat = 16'b1010011010000111 ;  
    10'd898     : sin_dat = 16'b1010011100010111 ;  
    10'd899     : sin_dat = 16'b1010011110100111 ;  
    10'd900     : sin_dat = 16'b1010100000111000 ;  
    10'd901     : sin_dat = 16'b1010100011001010 ;  
    10'd902     : sin_dat = 16'b1010100101011101 ;  
    10'd903     : sin_dat = 16'b1010100111110001 ;  
    10'd904     : sin_dat = 16'b1010101010000110 ;  
    10'd905     : sin_dat = 16'b1010101100011011 ;  
    10'd906     : sin_dat = 16'b1010101110110001 ;  
    10'd907     : sin_dat = 16'b1010110001001000 ;  
    10'd908     : sin_dat = 16'b1010110011100000 ;  
    10'd909     : sin_dat = 16'b1010110101111001 ;  
    10'd910     : sin_dat = 16'b1010111000010010 ;  
    10'd911     : sin_dat = 16'b1010111010101100 ;  
    10'd912     : sin_dat = 16'b1010111101000111 ;  
    10'd913     : sin_dat = 16'b1010111111100011 ;  
    10'd914     : sin_dat = 16'b1011000010000000 ;  
    10'd915     : sin_dat = 16'b1011000100011101 ;  
    10'd916     : sin_dat = 16'b1011000110111011 ;  
    10'd917     : sin_dat = 16'b1011001001011010 ;  
    10'd918     : sin_dat = 16'b1011001011111010 ;  
    10'd919     : sin_dat = 16'b1011001110011010 ;  
    10'd920     : sin_dat = 16'b1011010000111011 ;  
    10'd921     : sin_dat = 16'b1011010011011101 ;  
    10'd922     : sin_dat = 16'b1011010101111111 ;  
    10'd923     : sin_dat = 16'b1011011000100011 ;  
    10'd924     : sin_dat = 16'b1011011011000111 ;  
    10'd925     : sin_dat = 16'b1011011101101011 ;  
    10'd926     : sin_dat = 16'b1011100000010001 ;  
    10'd927     : sin_dat = 16'b1011100010110111 ;  
    10'd928     : sin_dat = 16'b1011100101011101 ;  
    10'd929     : sin_dat = 16'b1011101000000101 ;  
    10'd930     : sin_dat = 16'b1011101010101101 ;  
    10'd931     : sin_dat = 16'b1011101101010110 ;  
    10'd932     : sin_dat = 16'b1011101111111111 ;  
    10'd933     : sin_dat = 16'b1011110010101001 ;  
    10'd934     : sin_dat = 16'b1011110101010100 ;  
    10'd935     : sin_dat = 16'b1011110111111111 ;  
    10'd936     : sin_dat = 16'b1011111010101011 ;  
    10'd937     : sin_dat = 16'b1011111101011000 ;  
    10'd938     : sin_dat = 16'b1100000000000101 ;  
    10'd939     : sin_dat = 16'b1100000010110011 ;  
    10'd940     : sin_dat = 16'b1100000101100010 ;  
    10'd941     : sin_dat = 16'b1100001000010001 ;  
    10'd942     : sin_dat = 16'b1100001011000001 ;  
    10'd943     : sin_dat = 16'b1100001101110001 ;  
    10'd944     : sin_dat = 16'b1100010000100010 ;  
    10'd945     : sin_dat = 16'b1100010011010011 ;  
    10'd946     : sin_dat = 16'b1100010110000101 ;  
    10'd947     : sin_dat = 16'b1100011000111000 ;  
    10'd948     : sin_dat = 16'b1100011011101011 ;  
    10'd949     : sin_dat = 16'b1100011110011111 ;  
    10'd950     : sin_dat = 16'b1100100001010011 ;  
    10'd951     : sin_dat = 16'b1100100100001000 ;  
    10'd952     : sin_dat = 16'b1100100110111101 ;  
    10'd953     : sin_dat = 16'b1100101001110011 ;  
    10'd954     : sin_dat = 16'b1100101100101001 ;  
    10'd955     : sin_dat = 16'b1100101111100000 ;  
    10'd956     : sin_dat = 16'b1100110010010111 ;  
    10'd957     : sin_dat = 16'b1100110101001111 ;  
    10'd958     : sin_dat = 16'b1100111000001000 ;  
    10'd959     : sin_dat = 16'b1100111011000001 ;  
    10'd960     : sin_dat = 16'b1100111101111010 ;  
    10'd961     : sin_dat = 16'b1101000000110100 ;  
    10'd962     : sin_dat = 16'b1101000011101110 ;  
    10'd963     : sin_dat = 16'b1101000110101001 ;  
    10'd964     : sin_dat = 16'b1101001001100100 ;  
    10'd965     : sin_dat = 16'b1101001100011111 ;  
    10'd966     : sin_dat = 16'b1101001111011011 ;  
    10'd967     : sin_dat = 16'b1101010010011000 ;  
    10'd968     : sin_dat = 16'b1101010101010101 ;  
    10'd969     : sin_dat = 16'b1101011000010010 ;  
    10'd970     : sin_dat = 16'b1101011011010000 ;  
    10'd971     : sin_dat = 16'b1101011110001110 ;  
    10'd972     : sin_dat = 16'b1101100001001100 ;  
    10'd973     : sin_dat = 16'b1101100100001011 ;  
    10'd974     : sin_dat = 16'b1101100111001010 ;  
    10'd975     : sin_dat = 16'b1101101010001010 ;  
    10'd976     : sin_dat = 16'b1101101101001010 ;  
    10'd977     : sin_dat = 16'b1101110000001010 ;  
    10'd978     : sin_dat = 16'b1101110011001011 ;  
    10'd979     : sin_dat = 16'b1101110110001100 ;  
    10'd980     : sin_dat = 16'b1101111001001101 ;  
    10'd981     : sin_dat = 16'b1101111100001111 ;  
    10'd982     : sin_dat = 16'b1101111111010001 ;  
    10'd983     : sin_dat = 16'b1110000010010011 ;  
    10'd984     : sin_dat = 16'b1110000101010101 ;  
    10'd985     : sin_dat = 16'b1110001000011000 ;  
    10'd986     : sin_dat = 16'b1110001011011011 ;  
    10'd987     : sin_dat = 16'b1110001110011111 ;  
    10'd988     : sin_dat = 16'b1110010001100011 ;  
    10'd989     : sin_dat = 16'b1110010100100111 ;  
    10'd990     : sin_dat = 16'b1110010111101011 ;  
    10'd991     : sin_dat = 16'b1110011010101111 ;  
    10'd992     : sin_dat = 16'b1110011101110100 ;  
    10'd993     : sin_dat = 16'b1110100000111001 ;  
    10'd994     : sin_dat = 16'b1110100011111110 ;  
    10'd995     : sin_dat = 16'b1110100111000100 ;  
    10'd996     : sin_dat = 16'b1110101010001001 ;  
    10'd997     : sin_dat = 16'b1110101101001111 ;  
    10'd998     : sin_dat = 16'b1110110000010101 ;  
    10'd999     : sin_dat = 16'b1110110011011011 ;  
    10'd1000    : sin_dat = 16'b1110110110100010 ;  
    10'd1001    : sin_dat = 16'b1110111001101000 ;  
    10'd1002    : sin_dat = 16'b1110111100101111 ;  
    10'd1003    : sin_dat = 16'b1110111111110110 ;  
    10'd1004    : sin_dat = 16'b1111000010111101 ;  
    10'd1005    : sin_dat = 16'b1111000110000101 ;  
    10'd1006    : sin_dat = 16'b1111001001001100 ;  
    10'd1007    : sin_dat = 16'b1111001100010011 ;  
    10'd1008    : sin_dat = 16'b1111001111011011 ;  
    10'd1009    : sin_dat = 16'b1111010010100011 ;  
    10'd1010    : sin_dat = 16'b1111010101101011 ;  
    10'd1011    : sin_dat = 16'b1111011000110011 ;  
    10'd1012    : sin_dat = 16'b1111011011111011 ;  
    10'd1013    : sin_dat = 16'b1111011111000011 ;  
    10'd1014    : sin_dat = 16'b1111100010001011 ;  
    10'd1015    : sin_dat = 16'b1111100101010011 ;  
    10'd1016    : sin_dat = 16'b1111101000011100 ;  
    10'd1017    : sin_dat = 16'b1111101011100100 ;  
    10'd1018    : sin_dat = 16'b1111101110101101 ;  
    10'd1019    : sin_dat = 16'b1111110001110101 ;  
    10'd1020    : sin_dat = 16'b1111110100111110 ;  
    10'd1021    : sin_dat = 16'b1111111000000110 ;  
    10'd1022    : sin_dat = 16'b1111111011001111 ;  
    10'd1023    : sin_dat = 16'b1111111110010111 ;  
    default     : sin_dat = 16'd0;  
    endcase
end



//*******************************************************************************
//
// END of Module
//
//*******************************************************************************
endmodule
